VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_Burrows_Katie
  CLASS BLOCK ;
  FOREIGN tt_um_Burrows_Katie ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNADIFFAREA 17.639999 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
        RECT 156.550 -0.010 157.150 0.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 4.410000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
        RECT 134.470 -0.010 135.070 0.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 4.410000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
        RECT 112.390 -0.010 112.990 0.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 6.095000 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
        RECT 90.310 -0.010 90.910 0.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNAGATEAREA 4.000000 ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
        RECT 68.230 -0.010 68.830 0.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
        RECT 46.150 -0.010 46.750 0.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
        RECT 24.070 -0.010 24.670 0.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
        RECT 1.990 -0.010 2.590 0.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER pwell ;
        RECT 52.405 209.300 53.075 209.380 ;
        RECT 52.405 206.510 58.345 209.300 ;
      LAYER nwell ;
        RECT 97.880 207.490 104.300 212.770 ;
        RECT 105.960 207.490 112.380 212.770 ;
      LAYER pwell ;
        RECT 52.405 206.430 53.075 206.510 ;
        RECT 52.405 204.600 53.075 204.680 ;
        RECT 52.405 201.810 58.345 204.600 ;
      LAYER nwell ;
        RECT 63.065 203.420 65.485 206.700 ;
        RECT 92.045 203.455 94.465 206.735 ;
      LAYER pwell ;
        RECT 52.405 201.730 53.075 201.810 ;
      LAYER nwell ;
        RECT 97.880 200.500 104.300 205.780 ;
        RECT 105.960 200.500 112.380 205.780 ;
      LAYER pwell ;
        RECT 52.405 198.065 53.075 198.145 ;
        RECT 52.405 195.275 58.345 198.065 ;
        RECT 52.405 195.195 53.075 195.275 ;
      LAYER nwell ;
        RECT 76.590 194.110 83.010 199.390 ;
        RECT 97.880 193.510 104.300 198.790 ;
        RECT 105.960 193.510 112.380 198.790 ;
      LAYER pwell ;
        RECT 52.405 193.255 53.075 193.335 ;
        RECT 52.405 190.465 58.345 193.255 ;
        RECT 52.405 190.385 53.075 190.465 ;
      LAYER nwell ;
        RECT 76.590 187.195 83.010 192.475 ;
        RECT 97.880 186.485 104.300 191.765 ;
        RECT 105.960 186.485 112.380 191.765 ;
      LAYER pwell ;
        RECT 45.310 184.860 45.980 184.940 ;
        RECT 45.310 182.070 53.250 184.860 ;
        RECT 45.310 181.990 45.980 182.070 ;
        RECT 45.310 180.385 45.980 180.465 ;
        RECT 45.310 177.595 53.250 180.385 ;
        RECT 45.310 177.515 45.980 177.595 ;
        RECT 45.310 175.770 45.980 175.850 ;
        RECT 45.310 172.980 53.250 175.770 ;
        RECT 45.310 172.900 45.980 172.980 ;
        RECT 45.290 170.195 45.960 170.275 ;
        RECT 45.290 167.405 53.230 170.195 ;
      LAYER nwell ;
        RECT 88.440 169.485 90.860 172.765 ;
        RECT 106.185 167.870 112.605 173.150 ;
      LAYER pwell ;
        RECT 45.290 167.325 45.960 167.405 ;
        RECT 45.290 165.680 45.960 165.760 ;
        RECT 45.290 162.890 53.230 165.680 ;
        RECT 45.290 162.810 45.960 162.890 ;
        RECT 45.290 161.090 45.960 161.170 ;
        RECT 45.290 158.300 53.230 161.090 ;
      LAYER nwell ;
        RECT 88.435 159.485 90.855 162.765 ;
        RECT 106.185 160.760 112.605 166.040 ;
      LAYER pwell ;
        RECT 45.290 158.220 45.960 158.300 ;
        RECT 45.240 108.390 45.910 108.470 ;
        RECT 45.240 103.600 51.180 108.390 ;
        RECT 45.240 103.520 45.910 103.600 ;
      LAYER nwell ;
        RECT 54.505 103.410 60.925 108.690 ;
        RECT 64.655 103.410 71.075 108.690 ;
        RECT 73.935 103.365 80.355 108.645 ;
      LAYER pwell ;
        RECT 45.240 98.575 45.910 98.655 ;
        RECT 45.240 93.785 51.180 98.575 ;
        RECT 45.240 93.705 45.910 93.785 ;
      LAYER nwell ;
        RECT 54.505 93.515 60.925 98.795 ;
        RECT 64.655 93.535 71.075 98.815 ;
        RECT 73.935 93.475 80.355 98.755 ;
      LAYER pwell ;
        RECT 45.240 88.415 45.910 88.495 ;
        RECT 45.240 83.625 51.180 88.415 ;
        RECT 45.240 83.545 45.910 83.625 ;
      LAYER nwell ;
        RECT 54.505 83.470 60.925 88.750 ;
        RECT 64.655 83.595 71.075 88.875 ;
        RECT 73.890 83.640 80.310 88.920 ;
        RECT 97.335 82.380 103.755 95.350 ;
        RECT 115.680 82.380 122.100 95.350 ;
      LAYER pwell ;
        RECT 45.240 79.350 45.910 79.430 ;
        RECT 45.240 74.560 51.180 79.350 ;
        RECT 45.240 74.480 45.910 74.560 ;
      LAYER nwell ;
        RECT 54.505 74.270 60.925 79.550 ;
        RECT 64.655 74.175 71.075 79.455 ;
        RECT 73.935 74.080 80.355 79.360 ;
      LAYER pwell ;
        RECT 50.925 71.135 51.595 71.215 ;
        RECT 50.925 67.345 57.865 71.135 ;
        RECT 50.925 67.265 51.595 67.345 ;
        RECT 50.925 64.445 51.595 64.525 ;
        RECT 50.925 60.655 57.865 64.445 ;
        RECT 50.925 60.575 51.595 60.655 ;
        RECT 50.925 57.755 51.595 57.835 ;
        RECT 50.925 53.965 57.865 57.755 ;
      LAYER nwell ;
        RECT 63.850 55.615 72.270 69.355 ;
        RECT 76.205 56.035 84.625 69.835 ;
        RECT 97.030 64.090 103.450 77.060 ;
        RECT 115.685 63.845 122.105 76.815 ;
      LAYER pwell ;
        RECT 50.925 53.885 51.595 53.965 ;
        RECT 50.925 51.115 51.595 51.195 ;
        RECT 50.925 47.325 57.865 51.115 ;
        RECT 50.925 47.245 51.595 47.325 ;
        RECT 37.455 44.915 38.125 44.995 ;
        RECT 47.580 44.915 48.250 44.995 ;
        RECT 37.455 41.125 44.495 44.915 ;
        RECT 47.580 41.125 54.620 44.915 ;
        RECT 37.455 41.045 38.125 41.125 ;
        RECT 47.580 41.045 48.250 41.125 ;
      LAYER nwell ;
        RECT 64.105 38.910 72.525 52.650 ;
        RECT 76.225 38.390 84.645 52.190 ;
        RECT 112.870 44.815 121.290 57.155 ;
      LAYER pwell ;
        RECT 37.455 38.220 38.125 38.300 ;
        RECT 47.580 38.220 48.250 38.300 ;
        RECT 37.455 34.430 44.495 38.220 ;
        RECT 47.580 34.430 54.620 38.220 ;
        RECT 71.935 35.460 72.605 35.540 ;
        RECT 58.485 35.285 59.155 35.365 ;
        RECT 37.455 34.350 38.125 34.430 ;
        RECT 47.580 34.350 48.250 34.430 ;
        RECT 58.485 33.865 66.425 35.285 ;
        RECT 71.935 34.040 79.875 35.460 ;
        RECT 71.935 33.960 72.605 34.040 ;
        RECT 58.485 33.785 59.155 33.865 ;
        RECT 37.455 32.105 38.125 32.185 ;
        RECT 47.580 32.105 48.250 32.185 ;
        RECT 37.455 28.315 44.495 32.105 ;
        RECT 47.580 28.315 54.620 32.105 ;
        RECT 37.455 28.235 38.125 28.315 ;
        RECT 47.580 28.235 48.250 28.315 ;
        RECT 37.455 25.700 38.125 25.780 ;
        RECT 47.580 25.700 48.250 25.780 ;
        RECT 37.455 21.910 44.495 25.700 ;
        RECT 47.580 21.910 54.620 25.700 ;
        RECT 37.455 21.830 38.125 21.910 ;
        RECT 47.580 21.830 48.250 21.910 ;
      LAYER li1 ;
        RECT 98.755 212.750 99.285 213.280 ;
        RECT 107.035 212.750 107.565 213.280 ;
        RECT 98.870 212.355 99.170 212.750 ;
        RECT 98.565 212.185 103.315 212.355 ;
        RECT 103.750 211.690 104.080 212.435 ;
        RECT 107.150 212.355 107.450 212.750 ;
        RECT 106.645 212.185 111.395 212.355 ;
        RECT 104.365 211.690 104.895 211.825 ;
        RECT 103.750 211.360 104.895 211.690 ;
        RECT 52.575 208.385 52.905 209.210 ;
        RECT 53.610 209.130 54.310 210.320 ;
        RECT 97.360 210.090 97.960 210.690 ;
        RECT 53.340 208.960 58.090 209.130 ;
        RECT 51.665 207.685 52.905 208.385 ;
        RECT 52.575 206.600 52.905 207.685 ;
        RECT 58.770 207.540 59.300 208.070 ;
        RECT 98.565 207.905 103.315 208.075 ;
        RECT 103.000 207.490 103.170 207.905 ;
        RECT 103.750 207.825 104.080 211.360 ;
        RECT 104.365 211.295 104.895 211.360 ;
        RECT 111.830 211.535 112.160 212.435 ;
        RECT 112.465 211.535 112.995 211.675 ;
        RECT 111.830 211.205 112.995 211.535 ;
        RECT 105.555 210.230 106.155 210.830 ;
        RECT 106.645 207.905 111.395 208.075 ;
        RECT 106.850 207.760 107.155 207.905 ;
        RECT 111.830 207.825 112.160 211.205 ;
        RECT 112.465 211.145 112.995 211.205 ;
        RECT 106.855 207.490 107.155 207.760 ;
        RECT 53.340 206.680 58.090 206.850 ;
        RECT 63.870 206.750 64.400 207.280 ;
        RECT 92.955 206.750 93.485 207.280 ;
        RECT 102.820 206.960 103.350 207.490 ;
        RECT 106.740 206.960 107.270 207.490 ;
        RECT 53.410 206.350 53.710 206.680 ;
        RECT 53.295 205.820 53.825 206.350 ;
        RECT 63.985 206.285 64.155 206.750 ;
        RECT 64.955 206.365 65.285 206.385 ;
        RECT 63.790 206.115 64.460 206.285 ;
        RECT 52.575 203.485 52.905 204.510 ;
        RECT 53.600 204.430 54.300 205.255 ;
        RECT 62.330 205.040 63.220 205.930 ;
        RECT 53.340 204.260 58.090 204.430 ;
        RECT 63.790 203.940 64.460 204.005 ;
        RECT 51.665 202.785 52.905 203.485 ;
        RECT 63.775 203.835 64.460 203.940 ;
        RECT 63.775 203.475 64.175 203.835 ;
        RECT 64.935 203.755 65.285 206.365 ;
        RECT 93.080 206.320 93.380 206.750 ;
        RECT 92.770 206.150 93.440 206.320 ;
        RECT 93.080 206.115 93.380 206.150 ;
        RECT 91.240 205.040 92.130 205.930 ;
        RECT 92.770 203.870 93.440 204.040 ;
        RECT 93.915 203.930 94.245 206.400 ;
        RECT 98.755 205.555 99.285 206.085 ;
        RECT 107.035 205.555 107.565 206.085 ;
        RECT 98.870 205.365 99.170 205.555 ;
        RECT 98.565 205.195 103.315 205.365 ;
        RECT 58.770 202.885 59.300 203.415 ;
        RECT 63.690 202.945 64.220 203.475 ;
        RECT 52.575 201.900 52.905 202.785 ;
        RECT 64.955 202.400 65.285 203.755 ;
        RECT 93.080 203.495 93.380 203.870 ;
        RECT 93.890 203.790 94.245 203.930 ;
        RECT 103.750 204.770 104.080 205.445 ;
        RECT 107.150 205.365 107.450 205.555 ;
        RECT 106.645 205.195 111.395 205.365 ;
        RECT 104.385 204.770 104.915 204.910 ;
        RECT 103.750 204.440 104.915 204.770 ;
        RECT 92.955 202.965 93.485 203.495 ;
        RECT 93.890 202.495 94.220 203.790 ;
        RECT 97.360 202.915 97.960 203.515 ;
        RECT 53.340 201.980 58.090 202.150 ;
        RECT 53.370 201.540 53.670 201.980 ;
        RECT 64.955 201.970 65.495 202.400 ;
        RECT 64.965 201.870 65.495 201.970 ;
        RECT 93.765 201.965 94.295 202.495 ;
        RECT 53.255 201.010 53.785 201.540 ;
        RECT 98.565 200.915 103.315 201.085 ;
        RECT 103.085 200.425 103.255 200.915 ;
        RECT 103.750 200.835 104.080 204.440 ;
        RECT 104.385 204.380 104.915 204.440 ;
        RECT 111.830 204.770 112.160 205.445 ;
        RECT 112.465 204.770 112.995 204.910 ;
        RECT 111.830 204.440 112.995 204.770 ;
        RECT 105.555 203.150 106.155 203.750 ;
        RECT 106.645 200.915 111.395 201.085 ;
        RECT 106.940 200.425 107.240 200.915 ;
        RECT 111.830 200.835 112.160 204.440 ;
        RECT 112.465 204.380 112.995 204.440 ;
        RECT 81.235 198.975 81.935 200.195 ;
        RECT 102.905 199.895 103.435 200.425 ;
        RECT 106.825 199.895 107.355 200.425 ;
        RECT 52.575 196.950 52.905 197.975 ;
        RECT 53.525 197.895 54.225 198.825 ;
        RECT 77.275 198.805 82.025 198.975 ;
        RECT 82.460 198.935 82.790 199.055 ;
        RECT 82.460 198.235 83.760 198.935 ;
        RECT 98.755 198.580 99.285 199.110 ;
        RECT 107.035 198.650 107.565 199.180 ;
        RECT 98.870 198.375 99.170 198.580 ;
        RECT 53.340 197.725 58.090 197.895 ;
        RECT 51.665 196.250 52.905 196.950 ;
        RECT 58.770 196.490 59.300 197.020 ;
        RECT 76.035 196.505 76.565 197.035 ;
        RECT 52.575 195.365 52.905 196.250 ;
        RECT 53.340 195.445 58.090 195.615 ;
        RECT 53.425 195.120 53.725 195.445 ;
        RECT 53.310 194.590 53.840 195.120 ;
        RECT 77.275 194.525 82.025 194.695 ;
        RECT 77.595 194.140 77.895 194.525 ;
        RECT 82.460 194.445 82.790 198.235 ;
        RECT 98.565 198.205 103.315 198.375 ;
        RECT 103.750 197.595 104.080 198.455 ;
        RECT 107.150 198.375 107.450 198.650 ;
        RECT 106.645 198.205 111.395 198.375 ;
        RECT 104.385 197.595 104.915 197.800 ;
        RECT 103.750 197.270 104.915 197.595 ;
        RECT 111.830 197.595 112.160 198.455 ;
        RECT 112.465 197.595 112.995 197.800 ;
        RECT 111.830 197.270 112.995 197.595 ;
        RECT 103.750 197.265 104.815 197.270 ;
        RECT 111.830 197.265 112.895 197.270 ;
        RECT 97.360 195.965 97.960 196.565 ;
        RECT 52.575 192.260 52.905 193.165 ;
        RECT 53.580 193.085 54.280 193.900 ;
        RECT 77.480 193.610 78.010 194.140 ;
        RECT 98.565 193.925 103.315 194.095 ;
        RECT 103.085 193.545 103.255 193.925 ;
        RECT 103.750 193.845 104.080 197.265 ;
        RECT 105.555 196.280 106.155 196.880 ;
        RECT 106.645 193.925 111.395 194.095 ;
        RECT 106.940 193.545 107.240 193.925 ;
        RECT 111.830 193.845 112.160 197.265 ;
        RECT 53.340 192.915 58.090 193.085 ;
        RECT 51.665 191.560 52.905 192.260 ;
        RECT 81.235 192.060 81.935 193.090 ;
        RECT 102.905 193.015 103.435 193.545 ;
        RECT 106.825 193.015 107.355 193.545 ;
        RECT 52.575 190.555 52.905 191.560 ;
        RECT 58.770 191.445 59.300 191.975 ;
        RECT 77.275 191.890 82.025 192.060 ;
        RECT 82.460 192.040 82.790 192.140 ;
        RECT 82.460 191.340 83.760 192.040 ;
        RECT 98.755 191.605 99.285 192.135 ;
        RECT 107.035 191.670 107.565 192.200 ;
        RECT 98.935 191.350 99.105 191.605 ;
        RECT 53.340 190.635 58.090 190.805 ;
        RECT 53.390 190.300 53.690 190.635 ;
        RECT 53.310 189.770 53.840 190.300 ;
        RECT 76.015 189.230 76.545 189.760 ;
        RECT 77.275 187.610 82.025 187.780 ;
        RECT 77.595 187.275 77.895 187.610 ;
        RECT 82.460 187.530 82.790 191.340 ;
        RECT 98.565 191.180 103.315 191.350 ;
        RECT 103.750 190.495 104.080 191.430 ;
        RECT 107.150 191.350 107.450 191.670 ;
        RECT 106.645 191.180 111.395 191.350 ;
        RECT 104.385 190.495 104.915 190.735 ;
        RECT 103.750 190.205 104.915 190.495 ;
        RECT 103.750 190.165 104.815 190.205 ;
        RECT 97.360 188.940 97.960 189.540 ;
        RECT 77.480 186.745 78.010 187.275 ;
        RECT 98.565 186.900 103.315 187.070 ;
        RECT 103.085 186.385 103.255 186.900 ;
        RECT 103.750 186.820 104.080 190.165 ;
        RECT 111.830 190.055 112.160 191.430 ;
        RECT 112.465 190.055 112.995 190.295 ;
        RECT 111.830 189.765 112.995 190.055 ;
        RECT 111.830 189.725 112.895 189.765 ;
        RECT 105.555 188.940 106.155 189.540 ;
        RECT 106.645 186.900 111.395 187.070 ;
        RECT 106.940 186.385 107.240 186.900 ;
        RECT 111.830 186.820 112.160 189.725 ;
        RECT 45.480 184.690 45.810 184.770 ;
        RECT 46.345 184.690 47.045 185.865 ;
        RECT 102.905 185.855 103.435 186.385 ;
        RECT 106.825 185.855 107.355 186.385 ;
        RECT 44.420 183.990 45.810 184.690 ;
        RECT 46.225 184.520 53.015 184.690 ;
        RECT 45.480 182.160 45.810 183.990 ;
        RECT 53.630 183.175 54.160 183.705 ;
        RECT 46.225 182.240 53.015 182.410 ;
        RECT 52.710 181.880 53.010 182.240 ;
        RECT 52.620 181.350 53.150 181.880 ;
        RECT 58.315 181.160 58.485 183.040 ;
        RECT 118.650 182.370 118.820 183.040 ;
        RECT 45.480 180.235 45.810 180.295 ;
        RECT 44.420 179.535 45.810 180.235 ;
        RECT 46.345 180.215 47.045 181.135 ;
        RECT 46.225 180.045 53.015 180.215 ;
        RECT 45.480 177.685 45.810 179.535 ;
        RECT 53.630 178.720 54.160 179.250 ;
        RECT 58.315 178.740 58.485 180.620 ;
        RECT 118.650 179.950 118.820 181.830 ;
        RECT 46.225 177.765 53.015 177.935 ;
        RECT 52.705 177.365 53.005 177.765 ;
        RECT 52.620 176.835 53.150 177.365 ;
        RECT 45.480 175.635 45.810 175.680 ;
        RECT 44.420 174.935 45.810 175.635 ;
        RECT 46.345 175.600 47.045 176.570 ;
        RECT 58.315 176.320 58.485 178.200 ;
        RECT 118.650 177.530 118.820 179.410 ;
        RECT 118.650 176.320 118.820 176.990 ;
        RECT 46.225 175.430 53.015 175.600 ;
        RECT 45.480 173.070 45.810 174.935 ;
        RECT 53.630 174.025 54.160 174.555 ;
        RECT 46.225 173.150 53.015 173.320 ;
        RECT 52.710 172.765 53.010 173.150 ;
        RECT 52.620 172.235 53.150 172.765 ;
        RECT 89.020 172.735 89.550 173.265 ;
        RECT 106.770 172.735 107.470 173.755 ;
        RECT 89.165 172.350 89.465 172.735 ;
        RECT 106.770 172.630 111.620 172.735 ;
        RECT 106.870 172.565 111.620 172.630 ;
        RECT 89.165 172.180 89.835 172.350 ;
        RECT 89.165 172.120 89.465 172.180 ;
        RECT 45.460 170.090 45.790 170.105 ;
        RECT 44.420 169.390 45.790 170.090 ;
        RECT 46.260 170.025 46.960 171.000 ;
        RECT 87.665 170.730 88.555 171.620 ;
        RECT 90.310 171.375 90.640 172.430 ;
        RECT 112.055 172.075 112.385 172.815 ;
        RECT 112.055 171.375 113.500 172.075 ;
        RECT 90.310 170.675 91.575 171.375 ;
        RECT 46.205 169.855 52.995 170.025 ;
        RECT 89.165 169.900 89.835 170.070 ;
        RECT 45.460 167.495 45.790 169.390 ;
        RECT 89.165 169.295 89.465 169.900 ;
        RECT 90.310 169.820 90.640 170.675 ;
        RECT 105.525 169.875 106.125 170.475 ;
        RECT 53.605 168.315 54.135 168.845 ;
        RECT 89.045 168.765 89.575 169.295 ;
        RECT 106.970 168.455 107.670 168.465 ;
        RECT 106.870 168.285 111.620 168.455 ;
        RECT 46.205 167.575 52.995 167.745 ;
        RECT 45.460 165.450 45.790 165.590 ;
        RECT 46.260 165.510 46.960 166.550 ;
        RECT 52.275 166.540 52.975 167.575 ;
        RECT 106.970 167.340 107.670 168.285 ;
        RECT 112.055 168.205 112.385 171.375 ;
        RECT 106.770 165.625 107.470 166.585 ;
        RECT 106.770 165.535 111.620 165.625 ;
        RECT 44.485 164.750 45.790 165.450 ;
        RECT 46.205 165.340 52.995 165.510 ;
        RECT 106.870 165.455 111.620 165.535 ;
        RECT 112.055 165.520 112.385 165.705 ;
        RECT 45.460 162.980 45.790 164.750 ;
        RECT 112.055 164.820 113.410 165.520 ;
        RECT 53.635 164.005 54.165 164.535 ;
        RECT 46.205 163.060 52.995 163.230 ;
        RECT 52.275 162.000 52.975 163.060 ;
        RECT 89.035 162.675 89.565 163.205 ;
        RECT 93.760 162.705 94.290 163.235 ;
        RECT 105.525 163.085 106.125 163.685 ;
        RECT 89.170 162.350 89.470 162.675 ;
        RECT 89.160 162.180 89.830 162.350 ;
        RECT 89.170 162.110 89.470 162.180 ;
        RECT 45.460 160.985 45.790 161.000 ;
        RECT 44.420 160.285 45.790 160.985 ;
        RECT 46.260 160.920 46.960 161.975 ;
        RECT 46.205 160.750 52.995 160.920 ;
        RECT 87.755 160.770 88.645 161.660 ;
        RECT 90.305 161.420 90.635 162.430 ;
        RECT 45.460 158.390 45.790 160.285 ;
        RECT 90.305 160.720 91.640 161.420 ;
        RECT 106.870 161.175 111.620 161.345 ;
        RECT 53.615 159.405 54.145 159.935 ;
        RECT 89.160 159.900 89.830 160.070 ;
        RECT 89.170 159.305 89.470 159.900 ;
        RECT 90.305 159.820 90.635 160.720 ;
        RECT 106.970 160.200 107.670 161.175 ;
        RECT 112.055 161.095 112.385 164.820 ;
        RECT 89.045 158.775 89.575 159.305 ;
        RECT 46.205 158.470 52.995 158.640 ;
        RECT 52.255 157.250 52.955 158.470 ;
        RECT 45.675 153.500 45.845 155.380 ;
        RECT 110.680 154.710 110.850 155.380 ;
        RECT 45.675 151.080 45.845 152.960 ;
        RECT 110.680 152.290 110.850 154.170 ;
        RECT 45.675 148.660 45.845 150.540 ;
        RECT 110.680 149.870 110.850 151.750 ;
        RECT 45.675 146.240 45.845 148.120 ;
        RECT 110.680 147.450 110.850 149.330 ;
        RECT 45.675 143.820 45.845 145.700 ;
        RECT 110.680 145.030 110.850 146.910 ;
        RECT 45.675 141.400 45.845 143.280 ;
        RECT 110.680 142.610 110.850 144.490 ;
        RECT 45.675 138.980 45.845 140.860 ;
        RECT 110.680 140.190 110.850 142.070 ;
        RECT 45.675 136.560 45.845 138.440 ;
        RECT 110.680 137.770 110.850 139.650 ;
        RECT 110.680 136.560 110.850 137.230 ;
        RECT 46.045 108.900 46.575 109.070 ;
        RECT 55.030 108.910 55.560 109.080 ;
        RECT 65.265 108.910 65.795 109.080 ;
        RECT 45.410 107.055 45.740 108.300 ;
        RECT 46.220 108.220 46.390 108.900 ;
        RECT 55.205 108.275 55.375 108.910 ;
        RECT 46.175 108.050 50.925 108.220 ;
        RECT 55.190 108.105 59.940 108.275 ;
        RECT 46.220 108.045 46.390 108.050 ;
        RECT 44.055 106.055 45.740 107.055 ;
        RECT 60.375 106.480 60.705 108.355 ;
        RECT 65.440 108.275 65.610 108.910 ;
        RECT 65.340 108.105 70.090 108.275 ;
        RECT 70.525 106.520 70.855 108.355 ;
        RECT 78.655 108.230 79.355 109.660 ;
        RECT 74.620 108.060 79.370 108.230 ;
        RECT 78.655 108.050 79.355 108.060 ;
        RECT 45.410 103.690 45.740 106.055 ;
        RECT 51.585 105.915 52.115 106.445 ;
        RECT 60.375 106.410 61.750 106.480 ;
        RECT 70.525 106.410 71.960 106.520 ;
        RECT 60.375 106.240 62.035 106.410 ;
        RECT 70.525 106.240 72.060 106.410 ;
        RECT 60.375 106.150 61.750 106.240 ;
        RECT 70.525 106.190 71.960 106.240 ;
        RECT 54.025 103.950 54.555 104.480 ;
        RECT 46.175 103.770 50.925 103.940 ;
        RECT 55.190 103.825 59.940 103.995 ;
        RECT 46.245 103.320 46.415 103.770 ;
        RECT 55.230 103.355 55.400 103.825 ;
        RECT 60.375 103.745 60.705 106.150 ;
        RECT 64.185 103.920 64.715 104.450 ;
        RECT 65.340 103.825 70.090 103.995 ;
        RECT 45.785 102.320 46.785 103.320 ;
        RECT 54.770 102.355 55.770 103.355 ;
        RECT 65.725 103.295 65.895 103.825 ;
        RECT 70.525 103.745 70.855 106.190 ;
        RECT 73.385 105.710 73.915 106.240 ;
        RECT 74.620 103.780 79.370 103.950 ;
        RECT 65.265 102.295 66.265 103.295 ;
        RECT 74.640 103.275 74.810 103.780 ;
        RECT 74.235 102.385 75.125 103.275 ;
        RECT 79.805 102.740 80.135 108.310 ;
        RECT 82.960 104.415 83.130 105.085 ;
        RECT 79.520 102.695 80.135 102.740 ;
        RECT 79.420 102.525 80.135 102.695 ;
        RECT 79.520 102.410 80.135 102.525 ;
        RECT 82.960 101.995 83.130 103.875 ;
        RECT 123.795 103.205 123.965 105.085 ;
        RECT 46.045 100.050 46.575 100.220 ;
        RECT 45.410 97.260 45.740 98.485 ;
        RECT 46.220 98.405 46.390 100.050 ;
        RECT 55.030 98.950 55.560 99.120 ;
        RECT 65.265 98.970 65.795 99.140 ;
        RECT 46.175 98.235 50.925 98.405 ;
        RECT 55.205 98.380 55.375 98.950 ;
        RECT 55.190 98.210 59.940 98.380 ;
        RECT 44.055 96.260 45.740 97.260 ;
        RECT 45.410 93.875 45.740 96.260 ;
        RECT 51.605 95.805 52.135 96.335 ;
        RECT 60.375 96.090 60.705 98.460 ;
        RECT 65.440 98.400 65.610 98.970 ;
        RECT 64.185 97.725 64.715 98.255 ;
        RECT 65.340 98.230 70.090 98.400 ;
        RECT 70.525 96.195 70.855 98.480 ;
        RECT 78.655 98.340 79.355 99.755 ;
        RECT 82.960 99.575 83.130 101.455 ;
        RECT 123.795 100.785 123.965 102.665 ;
        RECT 123.795 99.575 123.965 100.245 ;
        RECT 74.620 98.170 79.370 98.340 ;
        RECT 78.655 98.145 79.355 98.170 ;
        RECT 60.375 96.060 61.795 96.090 ;
        RECT 70.525 96.060 71.960 96.195 ;
        RECT 60.375 95.890 62.035 96.060 ;
        RECT 70.525 95.890 72.060 96.060 ;
        RECT 60.375 95.760 61.795 95.890 ;
        RECT 70.525 95.865 71.960 95.890 ;
        RECT 46.175 93.955 50.925 94.125 ;
        RECT 54.025 94.020 54.555 94.550 ;
        RECT 46.245 93.410 46.415 93.955 ;
        RECT 55.190 93.930 59.940 94.100 ;
        RECT 55.230 93.445 55.400 93.930 ;
        RECT 60.375 93.850 60.705 95.760 ;
        RECT 65.340 93.950 70.090 94.120 ;
        RECT 45.785 92.410 46.785 93.410 ;
        RECT 54.770 92.445 55.770 93.445 ;
        RECT 65.725 93.400 65.895 93.950 ;
        RECT 70.525 93.870 70.855 95.865 ;
        RECT 73.405 95.745 73.935 96.275 ;
        RECT 74.620 93.890 79.370 94.060 ;
        RECT 65.265 92.400 66.265 93.400 ;
        RECT 74.640 93.375 74.810 93.890 ;
        RECT 74.235 92.485 75.125 93.375 ;
        RECT 79.805 93.225 80.135 98.420 ;
        RECT 93.250 95.685 93.780 96.215 ;
        RECT 96.455 95.620 97.455 96.620 ;
        RECT 112.285 96.280 112.815 96.810 ;
        RECT 98.145 95.840 98.675 96.010 ;
        RECT 94.550 93.920 95.550 94.895 ;
        RECT 96.215 94.735 96.745 94.760 ;
        RECT 96.215 94.590 96.830 94.735 ;
        RECT 96.585 94.565 96.830 94.590 ;
        RECT 94.550 93.895 96.390 93.920 ;
        RECT 95.125 93.750 96.390 93.895 ;
        RECT 79.520 93.175 80.135 93.225 ;
        RECT 79.420 93.005 80.135 93.175 ;
        RECT 79.520 92.895 80.135 93.005 ;
        RECT 93.520 92.330 94.520 93.330 ;
        RECT 96.220 93.260 96.390 93.750 ;
        RECT 96.660 93.675 96.830 94.565 ;
        RECT 97.180 94.295 97.350 95.620 ;
        RECT 98.325 94.935 98.495 95.840 ;
        RECT 114.785 95.620 115.785 96.620 ;
        RECT 116.475 95.840 117.005 96.010 ;
        RECT 98.020 94.765 102.770 94.935 ;
        RECT 98.020 94.295 102.770 94.305 ;
        RECT 97.180 94.135 102.770 94.295 ;
        RECT 97.180 94.125 98.150 94.135 ;
        RECT 103.205 93.770 103.535 95.015 ;
        RECT 104.585 93.770 105.585 94.210 ;
        RECT 112.880 93.920 113.880 94.895 ;
        RECT 114.545 94.735 115.075 94.760 ;
        RECT 114.545 94.590 115.160 94.735 ;
        RECT 114.915 94.565 115.160 94.590 ;
        RECT 112.880 93.895 114.720 93.920 ;
        RECT 96.660 93.505 102.770 93.675 ;
        RECT 103.205 93.440 105.585 93.770 ;
        RECT 113.455 93.750 114.720 93.895 ;
        RECT 96.220 93.090 97.720 93.260 ;
        RECT 95.165 92.920 95.780 93.090 ;
        RECT 95.610 92.855 95.780 92.920 ;
        RECT 97.550 93.045 97.720 93.090 ;
        RECT 97.550 92.875 102.770 93.045 ;
        RECT 95.610 92.685 97.260 92.855 ;
        RECT 97.090 92.615 97.260 92.685 ;
        RECT 97.090 92.445 97.735 92.615 ;
        RECT 94.350 92.225 94.520 92.330 ;
        RECT 97.565 92.415 97.735 92.445 ;
        RECT 97.565 92.245 102.770 92.415 ;
        RECT 94.350 92.055 97.155 92.225 ;
        RECT 91.170 90.825 92.170 91.825 ;
        RECT 96.985 91.785 97.155 92.055 ;
        RECT 93.410 91.575 96.795 91.745 ;
        RECT 96.985 91.615 102.770 91.785 ;
        RECT 93.410 91.510 93.580 91.575 ;
        RECT 93.050 91.340 93.580 91.510 ;
        RECT 94.205 91.050 96.070 91.220 ;
        RECT 89.850 90.610 90.380 90.695 ;
        RECT 89.850 90.440 90.640 90.610 ;
        RECT 90.470 90.040 90.640 90.440 ;
        RECT 91.820 90.500 91.990 90.825 ;
        RECT 94.205 90.500 94.375 91.050 ;
        RECT 91.820 90.330 94.375 90.500 ;
        RECT 95.900 90.525 96.070 91.050 ;
        RECT 96.625 91.155 96.795 91.575 ;
        RECT 96.625 90.985 102.770 91.155 ;
        RECT 95.900 90.355 102.770 90.525 ;
        RECT 91.460 90.040 93.735 90.065 ;
        RECT 55.030 89.180 55.560 89.350 ;
        RECT 65.265 89.305 65.795 89.475 ;
        RECT 46.045 88.830 46.575 89.000 ;
        RECT 45.410 87.900 45.740 88.325 ;
        RECT 46.220 88.245 46.390 88.830 ;
        RECT 55.215 88.335 55.385 89.180 ;
        RECT 65.450 88.460 65.620 89.305 ;
        RECT 46.175 88.075 50.925 88.245 ;
        RECT 55.190 88.165 59.940 88.335 ;
        RECT 44.055 86.900 45.740 87.900 ;
        RECT 45.410 83.715 45.740 86.900 ;
        RECT 51.585 85.730 52.115 86.260 ;
        RECT 60.375 86.105 60.705 88.415 ;
        RECT 65.340 88.290 70.090 88.460 ;
        RECT 64.185 87.720 64.715 88.250 ;
        RECT 70.525 86.255 70.855 88.540 ;
        RECT 78.605 88.505 79.305 89.945 ;
        RECT 90.470 89.895 93.735 90.040 ;
        RECT 90.470 89.870 91.630 89.895 ;
        RECT 93.565 89.725 102.770 89.895 ;
        RECT 87.955 89.265 88.955 89.665 ;
        RECT 87.955 89.095 102.770 89.265 ;
        RECT 87.955 88.665 88.955 89.095 ;
        RECT 98.020 88.605 102.770 88.635 ;
        RECT 74.575 88.335 79.325 88.505 ;
        RECT 70.525 86.200 71.960 86.255 ;
        RECT 60.375 86.040 61.840 86.105 ;
        RECT 60.375 85.870 62.035 86.040 ;
        RECT 70.525 86.030 72.060 86.200 ;
        RECT 70.525 85.925 71.960 86.030 ;
        RECT 73.345 85.985 73.875 86.515 ;
        RECT 60.375 85.775 61.840 85.870 ;
        RECT 54.025 83.970 54.555 84.500 ;
        RECT 46.175 83.795 50.925 83.965 ;
        RECT 55.190 83.885 59.940 84.055 ;
        RECT 46.245 83.255 46.415 83.795 ;
        RECT 55.230 83.430 55.400 83.885 ;
        RECT 60.375 83.805 60.705 85.775 ;
        RECT 65.340 84.010 70.090 84.180 ;
        RECT 65.725 83.545 65.895 84.010 ;
        RECT 70.525 83.930 70.855 85.925 ;
        RECT 74.575 84.055 79.325 84.225 ;
        RECT 74.580 83.695 74.750 84.055 ;
        RECT 45.785 82.255 46.785 83.255 ;
        RECT 54.770 82.430 55.770 83.430 ;
        RECT 65.265 82.545 66.265 83.545 ;
        RECT 74.310 82.695 75.310 83.695 ;
        RECT 79.760 82.820 80.090 88.585 ;
        RECT 96.480 88.465 102.770 88.605 ;
        RECT 96.480 88.435 98.235 88.465 ;
        RECT 96.480 88.335 96.650 88.435 ;
        RECT 89.850 88.165 96.650 88.335 ;
        RECT 97.045 88.005 98.185 88.020 ;
        RECT 97.045 87.850 102.770 88.005 ;
        RECT 97.045 87.800 97.215 87.850 ;
        RECT 98.020 87.835 102.770 87.850 ;
        RECT 90.905 87.630 97.215 87.800 ;
        RECT 90.905 87.285 91.075 87.630 ;
        RECT 98.020 87.355 102.770 87.375 ;
        RECT 97.505 87.315 102.770 87.355 ;
        RECT 90.490 86.285 91.490 87.285 ;
        RECT 92.630 87.205 102.770 87.315 ;
        RECT 92.630 87.185 98.175 87.205 ;
        RECT 92.630 87.145 97.675 87.185 ;
        RECT 92.630 86.870 92.800 87.145 ;
        RECT 92.185 86.700 92.800 86.870 ;
        RECT 93.285 86.575 102.770 86.745 ;
        RECT 93.285 85.860 93.455 86.575 ;
        RECT 94.750 85.945 102.770 86.115 ;
        RECT 92.565 84.860 93.565 85.860 ;
        RECT 94.750 85.350 94.920 85.945 ;
        RECT 94.290 85.180 94.920 85.350 ;
        RECT 94.470 85.140 94.920 85.180 ;
        RECT 95.460 85.315 102.770 85.485 ;
        RECT 95.460 84.445 95.630 85.315 ;
        RECT 93.440 84.275 95.630 84.445 ;
        RECT 96.070 84.685 102.770 84.855 ;
        RECT 93.440 83.915 93.610 84.275 ;
        RECT 92.565 83.330 93.610 83.915 ;
        RECT 96.070 83.595 96.240 84.685 ;
        RECT 94.675 83.525 96.240 83.595 ;
        RECT 94.495 83.425 96.240 83.525 ;
        RECT 96.690 84.055 102.770 84.225 ;
        RECT 94.495 83.355 95.025 83.425 ;
        RECT 92.565 82.915 93.565 83.330 ;
        RECT 96.690 83.040 96.860 84.055 ;
        RECT 79.385 82.655 80.090 82.820 ;
        RECT 95.630 82.870 96.860 83.040 ;
        RECT 97.180 83.425 102.770 83.595 ;
        RECT 79.385 82.650 79.915 82.655 ;
        RECT 95.630 82.375 95.800 82.870 ;
        RECT 94.835 81.375 95.835 82.375 ;
        RECT 97.180 82.100 97.350 83.425 ;
        RECT 98.020 82.795 102.770 82.965 ;
        RECT 98.405 82.375 98.575 82.795 ;
        RECT 103.205 82.715 103.535 93.440 ;
        RECT 104.585 93.210 105.585 93.440 ;
        RECT 111.850 92.330 112.850 93.330 ;
        RECT 114.550 93.260 114.720 93.750 ;
        RECT 114.990 93.675 115.160 94.565 ;
        RECT 115.510 94.295 115.680 95.620 ;
        RECT 116.655 94.935 116.825 95.840 ;
        RECT 116.365 94.765 121.115 94.935 ;
        RECT 116.365 94.295 121.115 94.305 ;
        RECT 115.510 94.135 121.115 94.295 ;
        RECT 115.510 94.125 116.480 94.135 ;
        RECT 114.990 93.505 121.115 93.675 ;
        RECT 114.550 93.090 116.050 93.260 ;
        RECT 113.495 92.920 114.110 93.090 ;
        RECT 113.940 92.855 114.110 92.920 ;
        RECT 115.880 93.045 116.050 93.090 ;
        RECT 115.880 92.875 121.115 93.045 ;
        RECT 113.940 92.685 115.590 92.855 ;
        RECT 115.420 92.615 115.590 92.685 ;
        RECT 115.420 92.445 116.065 92.615 ;
        RECT 112.680 92.225 112.850 92.330 ;
        RECT 115.895 92.415 116.065 92.445 ;
        RECT 115.895 92.245 121.115 92.415 ;
        RECT 112.680 92.055 115.485 92.225 ;
        RECT 109.500 90.825 110.500 91.825 ;
        RECT 115.315 91.785 115.485 92.055 ;
        RECT 111.740 91.575 115.125 91.745 ;
        RECT 115.315 91.615 121.115 91.785 ;
        RECT 111.740 91.510 111.910 91.575 ;
        RECT 111.380 91.340 111.910 91.510 ;
        RECT 112.535 91.050 114.400 91.220 ;
        RECT 108.180 90.610 108.710 90.695 ;
        RECT 108.180 90.440 108.970 90.610 ;
        RECT 108.800 90.040 108.970 90.440 ;
        RECT 110.150 90.500 110.320 90.825 ;
        RECT 112.535 90.500 112.705 91.050 ;
        RECT 110.150 90.330 112.705 90.500 ;
        RECT 114.230 90.525 114.400 91.050 ;
        RECT 114.955 91.155 115.125 91.575 ;
        RECT 114.955 90.985 121.115 91.155 ;
        RECT 114.230 90.355 121.115 90.525 ;
        RECT 109.790 90.040 112.065 90.065 ;
        RECT 108.800 89.895 112.065 90.040 ;
        RECT 108.800 89.870 109.960 89.895 ;
        RECT 111.895 89.725 121.115 89.895 ;
        RECT 106.285 89.265 107.285 89.685 ;
        RECT 121.550 89.640 121.880 95.015 ;
        RECT 106.285 89.095 121.115 89.265 ;
        RECT 106.285 88.685 107.285 89.095 ;
        RECT 121.550 88.940 122.995 89.640 ;
        RECT 116.365 88.605 121.115 88.635 ;
        RECT 114.810 88.465 121.115 88.605 ;
        RECT 114.810 88.435 116.565 88.465 ;
        RECT 114.810 88.335 114.980 88.435 ;
        RECT 108.180 88.165 114.980 88.335 ;
        RECT 115.375 88.005 116.515 88.020 ;
        RECT 115.375 87.850 121.115 88.005 ;
        RECT 115.375 87.800 115.545 87.850 ;
        RECT 116.365 87.835 121.115 87.850 ;
        RECT 109.235 87.630 115.545 87.800 ;
        RECT 109.235 87.285 109.405 87.630 ;
        RECT 116.365 87.355 121.115 87.375 ;
        RECT 115.835 87.315 121.115 87.355 ;
        RECT 108.820 86.285 109.820 87.285 ;
        RECT 110.960 87.205 121.115 87.315 ;
        RECT 110.960 87.185 116.505 87.205 ;
        RECT 110.960 87.145 116.005 87.185 ;
        RECT 110.960 86.870 111.130 87.145 ;
        RECT 110.515 86.700 111.130 86.870 ;
        RECT 111.615 86.575 121.115 86.745 ;
        RECT 111.615 85.860 111.785 86.575 ;
        RECT 113.080 85.945 121.115 86.115 ;
        RECT 110.895 84.860 111.895 85.860 ;
        RECT 113.080 85.350 113.250 85.945 ;
        RECT 112.620 85.180 113.250 85.350 ;
        RECT 112.800 85.140 113.250 85.180 ;
        RECT 113.790 85.315 121.115 85.485 ;
        RECT 113.790 84.445 113.960 85.315 ;
        RECT 111.770 84.275 113.960 84.445 ;
        RECT 114.400 84.685 121.115 84.855 ;
        RECT 111.770 83.915 111.940 84.275 ;
        RECT 110.895 83.330 111.940 83.915 ;
        RECT 114.400 83.595 114.570 84.685 ;
        RECT 113.005 83.525 114.570 83.595 ;
        RECT 112.825 83.425 114.570 83.525 ;
        RECT 115.020 84.055 121.115 84.225 ;
        RECT 112.825 83.355 113.355 83.425 ;
        RECT 110.895 82.915 111.895 83.330 ;
        RECT 115.020 83.040 115.190 84.055 ;
        RECT 113.960 82.870 115.190 83.040 ;
        RECT 115.510 83.425 121.115 83.595 ;
        RECT 113.960 82.375 114.130 82.870 ;
        RECT 96.755 82.065 97.350 82.100 ;
        RECT 96.575 81.930 97.350 82.065 ;
        RECT 96.575 81.895 97.105 81.930 ;
        RECT 97.990 81.375 98.990 82.375 ;
        RECT 113.165 81.375 114.165 82.375 ;
        RECT 115.510 82.100 115.680 83.425 ;
        RECT 116.365 82.795 121.115 82.965 ;
        RECT 116.735 82.375 116.905 82.795 ;
        RECT 121.550 82.715 121.880 88.940 ;
        RECT 115.085 82.065 115.680 82.100 ;
        RECT 114.905 81.930 115.680 82.065 ;
        RECT 114.905 81.895 115.435 81.930 ;
        RECT 116.320 81.375 117.320 82.375 ;
        RECT 46.045 79.755 46.575 79.925 ;
        RECT 45.410 77.330 45.740 79.260 ;
        RECT 46.220 79.180 46.390 79.755 ;
        RECT 55.030 79.745 55.560 79.915 ;
        RECT 65.265 79.790 65.795 79.960 ;
        RECT 46.175 79.010 50.925 79.180 ;
        RECT 55.205 79.135 55.375 79.745 ;
        RECT 54.025 78.550 54.555 79.080 ;
        RECT 55.190 78.965 59.940 79.135 ;
        RECT 43.685 76.330 45.740 77.330 ;
        RECT 60.375 77.155 60.705 79.215 ;
        RECT 65.440 79.040 65.610 79.790 ;
        RECT 78.855 79.645 79.385 79.650 ;
        RECT 78.675 79.480 79.385 79.645 ;
        RECT 64.185 78.455 64.715 78.985 ;
        RECT 65.340 78.870 70.090 79.040 ;
        RECT 60.375 77.105 61.805 77.155 ;
        RECT 51.605 76.530 52.135 77.060 ;
        RECT 60.375 76.935 62.035 77.105 ;
        RECT 60.375 76.825 61.805 76.935 ;
        RECT 70.525 76.925 70.855 79.120 ;
        RECT 78.675 78.945 79.375 79.480 ;
        RECT 74.620 78.775 79.375 78.945 ;
        RECT 78.675 78.760 79.375 78.775 ;
        RECT 70.525 76.875 71.735 76.925 ;
        RECT 45.410 74.650 45.740 76.330 ;
        RECT 46.175 74.730 50.925 74.900 ;
        RECT 46.245 74.250 46.415 74.730 ;
        RECT 55.190 74.685 59.940 74.855 ;
        RECT 45.785 73.250 46.785 74.250 ;
        RECT 55.230 74.225 55.400 74.685 ;
        RECT 60.375 74.605 60.705 76.825 ;
        RECT 70.525 76.705 72.060 76.875 ;
        RECT 70.525 76.595 71.735 76.705 ;
        RECT 65.340 74.590 70.090 74.760 ;
        RECT 65.725 74.370 65.895 74.590 ;
        RECT 70.525 74.510 70.855 76.595 ;
        RECT 73.365 76.285 73.895 76.815 ;
        RECT 74.630 74.665 74.800 74.685 ;
        RECT 74.620 74.495 79.370 74.665 ;
        RECT 54.770 73.225 55.770 74.225 ;
        RECT 65.265 73.370 66.265 74.370 ;
        RECT 74.630 74.070 74.800 74.495 ;
        RECT 73.905 73.070 74.905 74.070 ;
        RECT 79.805 73.380 80.135 79.025 ;
        RECT 92.940 77.300 93.470 77.830 ;
        RECT 96.215 77.330 97.215 78.330 ;
        RECT 97.855 77.550 98.385 77.720 ;
        RECT 94.260 75.630 95.260 76.605 ;
        RECT 95.925 76.445 96.455 76.470 ;
        RECT 95.925 76.300 96.540 76.445 ;
        RECT 96.295 76.275 96.540 76.300 ;
        RECT 94.260 75.605 96.100 75.630 ;
        RECT 94.835 75.460 96.100 75.605 ;
        RECT 93.230 74.040 94.230 75.040 ;
        RECT 95.930 74.970 96.100 75.460 ;
        RECT 96.370 75.385 96.540 76.275 ;
        RECT 96.890 76.005 97.060 77.330 ;
        RECT 98.035 76.645 98.205 77.550 ;
        RECT 111.590 76.925 112.120 77.455 ;
        RECT 114.815 77.085 115.815 78.085 ;
        RECT 116.505 77.305 117.035 77.475 ;
        RECT 97.715 76.475 102.465 76.645 ;
        RECT 97.715 76.005 102.465 76.015 ;
        RECT 96.890 75.845 102.465 76.005 ;
        RECT 96.890 75.835 97.860 75.845 ;
        RECT 96.370 75.215 102.465 75.385 ;
        RECT 95.930 74.800 97.430 74.970 ;
        RECT 94.875 74.630 95.490 74.800 ;
        RECT 95.320 74.565 95.490 74.630 ;
        RECT 97.260 74.755 97.430 74.800 ;
        RECT 97.260 74.585 102.465 74.755 ;
        RECT 95.320 74.395 96.970 74.565 ;
        RECT 96.800 74.325 96.970 74.395 ;
        RECT 96.800 74.155 97.445 74.325 ;
        RECT 94.060 73.935 94.230 74.040 ;
        RECT 97.275 74.125 97.445 74.155 ;
        RECT 97.275 73.955 102.465 74.125 ;
        RECT 94.060 73.765 96.865 73.935 ;
        RECT 79.515 73.050 80.135 73.380 ;
        RECT 90.880 72.535 91.880 73.535 ;
        RECT 96.695 73.495 96.865 73.765 ;
        RECT 93.120 73.285 96.505 73.455 ;
        RECT 96.695 73.325 102.465 73.495 ;
        RECT 93.120 73.220 93.290 73.285 ;
        RECT 92.760 73.050 93.290 73.220 ;
        RECT 93.915 72.760 95.780 72.930 ;
        RECT 89.560 72.320 90.090 72.405 ;
        RECT 89.560 72.150 90.350 72.320 ;
        RECT 51.095 71.920 52.160 72.015 ;
        RECT 51.095 71.750 52.260 71.920 ;
        RECT 90.180 71.750 90.350 72.150 ;
        RECT 91.530 72.210 91.700 72.535 ;
        RECT 93.915 72.210 94.085 72.760 ;
        RECT 91.530 72.040 94.085 72.210 ;
        RECT 95.610 72.235 95.780 72.760 ;
        RECT 96.335 72.865 96.505 73.285 ;
        RECT 96.335 72.695 102.465 72.865 ;
        RECT 95.610 72.065 102.465 72.235 ;
        RECT 91.170 71.750 93.445 71.775 ;
        RECT 51.095 71.685 52.160 71.750 ;
        RECT 51.095 67.435 51.425 71.685 ;
        RECT 51.860 70.965 52.030 71.685 ;
        RECT 90.180 71.605 93.445 71.750 ;
        RECT 90.180 71.580 91.340 71.605 ;
        RECT 93.275 71.435 102.465 71.605 ;
        RECT 87.665 70.975 88.665 71.395 ;
        RECT 51.850 70.795 57.620 70.965 ;
        RECT 87.665 70.805 102.465 70.975 ;
        RECT 87.665 70.395 88.665 70.805 ;
        RECT 97.715 70.315 102.465 70.345 ;
        RECT 96.190 70.175 102.465 70.315 ;
        RECT 96.190 70.145 97.945 70.175 ;
        RECT 96.190 70.045 96.360 70.145 ;
        RECT 89.560 69.875 96.360 70.045 ;
        RECT 96.755 69.715 97.895 69.730 ;
        RECT 75.650 69.420 76.180 69.595 ;
        RECT 96.755 69.560 102.465 69.715 ;
        RECT 96.755 69.510 96.925 69.560 ;
        RECT 97.715 69.545 102.465 69.560 ;
        RECT 75.650 69.250 83.660 69.420 ;
        RECT 75.650 69.065 76.180 69.250 ;
        RECT 63.905 68.950 64.635 68.955 ;
        RECT 63.725 68.940 64.635 68.950 ;
        RECT 58.260 68.275 58.790 68.805 ;
        RECT 63.725 68.785 71.305 68.940 ;
        RECT 63.725 68.780 64.255 68.785 ;
        RECT 64.515 68.770 71.305 68.785 ;
        RECT 61.575 67.860 71.305 68.030 ;
        RECT 51.850 67.665 57.620 67.685 ;
        RECT 51.840 67.515 57.620 67.665 ;
        RECT 51.840 67.050 52.010 67.515 ;
        RECT 51.380 66.050 52.380 67.050 ;
        RECT 61.575 66.210 61.745 67.860 ;
        RECT 63.905 67.130 64.765 67.135 ;
        RECT 63.725 67.120 64.765 67.130 ;
        RECT 63.725 66.965 71.305 67.120 ;
        RECT 63.725 66.960 64.255 66.965 ;
        RECT 64.515 66.950 71.305 66.965 ;
        RECT 61.575 66.040 71.305 66.210 ;
        RECT 51.095 65.380 52.160 65.410 ;
        RECT 51.095 65.210 52.260 65.380 ;
        RECT 51.095 65.080 52.160 65.210 ;
        RECT 51.095 60.745 51.425 65.080 ;
        RECT 51.850 64.275 52.020 65.080 ;
        RECT 61.575 64.390 61.745 66.040 ;
        RECT 63.905 65.310 64.745 65.315 ;
        RECT 63.725 65.300 64.745 65.310 ;
        RECT 63.725 65.145 71.305 65.300 ;
        RECT 63.725 65.140 64.255 65.145 ;
        RECT 64.515 65.130 71.305 65.145 ;
        RECT 51.850 64.105 57.620 64.275 ;
        RECT 61.575 64.220 71.305 64.390 ;
        RECT 58.280 62.940 58.810 63.470 ;
        RECT 61.575 62.570 61.745 64.220 ;
        RECT 63.735 63.480 64.635 63.495 ;
        RECT 63.735 63.325 71.305 63.480 ;
        RECT 64.515 63.310 71.305 63.325 ;
        RECT 61.575 62.400 71.305 62.570 ;
        RECT 51.850 60.975 57.620 60.995 ;
        RECT 51.840 60.825 57.620 60.975 ;
        RECT 51.840 60.360 52.010 60.825 ;
        RECT 61.575 60.750 61.745 62.400 ;
        RECT 63.735 61.660 64.265 61.670 ;
        RECT 63.735 61.500 71.305 61.660 ;
        RECT 63.915 61.490 71.305 61.500 ;
        RECT 61.575 60.580 71.305 60.750 ;
        RECT 51.380 59.360 52.380 60.360 ;
        RECT 61.575 58.930 61.745 60.580 ;
        RECT 63.915 59.845 64.780 59.855 ;
        RECT 63.735 59.840 64.780 59.845 ;
        RECT 63.735 59.685 71.305 59.840 ;
        RECT 63.735 59.675 64.265 59.685 ;
        RECT 64.515 59.670 71.305 59.685 ;
        RECT 61.575 58.760 71.305 58.930 ;
        RECT 51.095 58.685 52.160 58.755 ;
        RECT 51.095 58.515 52.260 58.685 ;
        RECT 51.095 58.425 52.160 58.515 ;
        RECT 51.095 54.055 51.425 58.425 ;
        RECT 51.855 57.585 52.025 58.425 ;
        RECT 61.575 57.920 61.745 58.760 ;
        RECT 63.725 58.020 64.770 58.035 ;
        RECT 62.145 57.920 62.415 58.005 ;
        RECT 61.575 57.750 62.415 57.920 ;
        RECT 63.725 57.865 71.305 58.020 ;
        RECT 64.515 57.850 71.305 57.865 ;
        RECT 51.850 57.415 57.620 57.585 ;
        RECT 61.575 57.110 61.745 57.750 ;
        RECT 62.145 57.675 62.415 57.750 ;
        RECT 61.575 56.940 71.305 57.110 ;
        RECT 61.575 56.210 61.745 56.940 ;
        RECT 64.000 56.215 64.195 56.330 ;
        RECT 64.000 56.210 64.730 56.215 ;
        RECT 61.430 56.040 61.960 56.210 ;
        RECT 63.735 56.200 64.730 56.210 ;
        RECT 63.735 56.045 71.305 56.200 ;
        RECT 71.720 56.185 72.050 69.020 ;
        RECT 74.450 67.970 83.660 68.140 ;
        RECT 74.500 65.580 74.670 67.970 ;
        RECT 75.650 66.860 76.180 67.080 ;
        RECT 75.650 66.690 83.660 66.860 ;
        RECT 75.650 66.550 76.180 66.690 ;
        RECT 74.500 65.410 83.660 65.580 ;
        RECT 74.500 63.020 74.670 65.410 ;
        RECT 75.650 64.300 76.180 64.475 ;
        RECT 75.650 64.130 83.660 64.300 ;
        RECT 75.650 63.945 76.180 64.130 ;
        RECT 74.500 62.850 83.660 63.020 ;
        RECT 74.500 60.460 74.670 62.850 ;
        RECT 75.650 61.740 76.180 61.945 ;
        RECT 75.650 61.570 83.660 61.740 ;
        RECT 75.650 61.415 76.180 61.570 ;
        RECT 74.500 60.290 83.660 60.460 ;
        RECT 74.500 57.900 74.670 60.290 ;
        RECT 75.650 59.180 76.180 59.300 ;
        RECT 75.650 59.010 83.660 59.180 ;
        RECT 75.650 58.770 76.180 59.010 ;
        RECT 74.500 57.730 83.660 57.900 ;
        RECT 74.500 57.320 74.670 57.730 ;
        RECT 74.500 57.170 74.775 57.320 ;
        RECT 74.505 56.990 74.775 57.170 ;
        RECT 63.735 56.040 64.265 56.045 ;
        RECT 64.515 56.030 71.305 56.045 ;
        RECT 71.700 55.950 72.050 56.185 ;
        RECT 74.530 56.155 74.700 56.990 ;
        RECT 75.650 56.620 76.180 56.825 ;
        RECT 75.650 56.450 83.660 56.620 ;
        RECT 75.650 56.295 76.180 56.450 ;
        RECT 84.075 56.370 84.405 69.500 ;
        RECT 90.615 69.340 96.925 69.510 ;
        RECT 90.615 68.995 90.785 69.340 ;
        RECT 97.715 69.065 102.465 69.085 ;
        RECT 97.215 69.025 102.465 69.065 ;
        RECT 90.200 67.995 91.200 68.995 ;
        RECT 92.340 68.915 102.465 69.025 ;
        RECT 92.340 68.895 97.885 68.915 ;
        RECT 92.340 68.855 97.385 68.895 ;
        RECT 92.340 68.580 92.510 68.855 ;
        RECT 91.895 68.410 92.510 68.580 ;
        RECT 92.995 68.285 102.465 68.455 ;
        RECT 92.995 67.570 93.165 68.285 ;
        RECT 94.460 67.655 102.465 67.825 ;
        RECT 92.275 66.570 93.275 67.570 ;
        RECT 94.460 67.060 94.630 67.655 ;
        RECT 94.000 66.890 94.630 67.060 ;
        RECT 94.180 66.850 94.630 66.890 ;
        RECT 95.170 67.025 102.465 67.195 ;
        RECT 95.170 66.155 95.340 67.025 ;
        RECT 93.150 65.985 95.340 66.155 ;
        RECT 95.780 66.395 102.465 66.565 ;
        RECT 93.150 65.625 93.320 65.985 ;
        RECT 92.275 65.040 93.320 65.625 ;
        RECT 95.780 65.305 95.950 66.395 ;
        RECT 94.385 65.235 95.950 65.305 ;
        RECT 94.205 65.135 95.950 65.235 ;
        RECT 96.400 65.765 102.465 65.935 ;
        RECT 94.205 65.065 94.735 65.135 ;
        RECT 92.275 64.625 93.275 65.040 ;
        RECT 96.400 64.750 96.570 65.765 ;
        RECT 102.900 65.480 103.230 76.725 ;
        RECT 112.910 75.385 113.910 76.360 ;
        RECT 114.575 76.200 115.105 76.225 ;
        RECT 114.575 76.055 115.190 76.200 ;
        RECT 114.945 76.030 115.190 76.055 ;
        RECT 112.910 75.360 114.750 75.385 ;
        RECT 113.485 75.215 114.750 75.360 ;
        RECT 111.880 73.795 112.880 74.795 ;
        RECT 114.580 74.725 114.750 75.215 ;
        RECT 115.020 75.140 115.190 76.030 ;
        RECT 115.540 75.760 115.710 77.085 ;
        RECT 116.685 76.400 116.855 77.305 ;
        RECT 116.370 76.230 121.120 76.400 ;
        RECT 116.370 75.760 121.120 75.770 ;
        RECT 115.540 75.600 121.120 75.760 ;
        RECT 115.540 75.590 116.510 75.600 ;
        RECT 115.020 74.970 121.120 75.140 ;
        RECT 114.580 74.555 116.080 74.725 ;
        RECT 113.525 74.385 114.140 74.555 ;
        RECT 113.970 74.320 114.140 74.385 ;
        RECT 115.910 74.510 116.080 74.555 ;
        RECT 115.910 74.340 121.120 74.510 ;
        RECT 113.970 74.150 115.620 74.320 ;
        RECT 115.450 74.080 115.620 74.150 ;
        RECT 115.450 73.910 116.095 74.080 ;
        RECT 112.710 73.690 112.880 73.795 ;
        RECT 115.925 73.880 116.095 73.910 ;
        RECT 115.925 73.710 121.120 73.880 ;
        RECT 112.710 73.520 115.515 73.690 ;
        RECT 109.530 72.290 110.530 73.290 ;
        RECT 115.345 73.250 115.515 73.520 ;
        RECT 111.770 73.040 115.155 73.210 ;
        RECT 115.345 73.080 121.120 73.250 ;
        RECT 111.770 72.975 111.940 73.040 ;
        RECT 111.410 72.805 111.940 72.975 ;
        RECT 112.565 72.515 114.430 72.685 ;
        RECT 108.210 72.075 108.740 72.160 ;
        RECT 108.210 71.905 109.000 72.075 ;
        RECT 108.830 71.505 109.000 71.905 ;
        RECT 110.180 71.965 110.350 72.290 ;
        RECT 112.565 71.965 112.735 72.515 ;
        RECT 110.180 71.795 112.735 71.965 ;
        RECT 114.260 71.990 114.430 72.515 ;
        RECT 114.985 72.620 115.155 73.040 ;
        RECT 114.985 72.450 121.120 72.620 ;
        RECT 114.260 71.820 121.120 71.990 ;
        RECT 109.820 71.505 112.095 71.530 ;
        RECT 108.830 71.360 112.095 71.505 ;
        RECT 108.830 71.335 109.990 71.360 ;
        RECT 111.925 71.190 121.120 71.360 ;
        RECT 106.315 70.730 107.315 71.165 ;
        RECT 121.555 71.035 121.885 76.480 ;
        RECT 106.315 70.560 121.120 70.730 ;
        RECT 106.315 70.165 107.315 70.560 ;
        RECT 121.555 70.335 122.720 71.035 ;
        RECT 116.370 70.070 121.120 70.100 ;
        RECT 114.840 69.930 121.120 70.070 ;
        RECT 114.840 69.900 116.595 69.930 ;
        RECT 114.840 69.800 115.010 69.900 ;
        RECT 108.210 69.630 115.010 69.800 ;
        RECT 115.405 69.470 116.545 69.485 ;
        RECT 115.405 69.315 121.120 69.470 ;
        RECT 115.405 69.265 115.575 69.315 ;
        RECT 116.370 69.300 121.120 69.315 ;
        RECT 109.265 69.095 115.575 69.265 ;
        RECT 109.265 68.750 109.435 69.095 ;
        RECT 116.370 68.820 121.120 68.840 ;
        RECT 115.865 68.780 121.120 68.820 ;
        RECT 108.850 67.750 109.850 68.750 ;
        RECT 110.990 68.670 121.120 68.780 ;
        RECT 110.990 68.650 116.535 68.670 ;
        RECT 110.990 68.610 116.035 68.650 ;
        RECT 110.990 68.335 111.160 68.610 ;
        RECT 110.545 68.165 111.160 68.335 ;
        RECT 111.645 68.040 121.120 68.210 ;
        RECT 111.645 67.325 111.815 68.040 ;
        RECT 113.110 67.410 121.120 67.580 ;
        RECT 110.925 66.325 111.925 67.325 ;
        RECT 113.110 66.815 113.280 67.410 ;
        RECT 112.650 66.645 113.280 66.815 ;
        RECT 112.830 66.605 113.280 66.645 ;
        RECT 113.820 66.780 121.120 66.950 ;
        RECT 113.820 65.910 113.990 66.780 ;
        RECT 111.800 65.740 113.990 65.910 ;
        RECT 114.430 66.150 121.120 66.320 ;
        RECT 104.090 65.480 104.620 65.595 ;
        RECT 95.340 64.580 96.570 64.750 ;
        RECT 96.890 65.135 102.465 65.305 ;
        RECT 102.900 65.180 104.620 65.480 ;
        RECT 111.800 65.380 111.970 65.740 ;
        RECT 95.340 64.085 95.510 64.580 ;
        RECT 94.545 63.085 95.545 64.085 ;
        RECT 96.890 63.810 97.060 65.135 ;
        RECT 97.715 64.505 102.465 64.675 ;
        RECT 98.115 64.085 98.285 64.505 ;
        RECT 102.900 64.425 103.230 65.180 ;
        RECT 104.090 65.065 104.620 65.180 ;
        RECT 110.925 64.795 111.970 65.380 ;
        RECT 114.430 65.060 114.600 66.150 ;
        RECT 113.035 64.990 114.600 65.060 ;
        RECT 112.855 64.890 114.600 64.990 ;
        RECT 115.050 65.520 121.120 65.690 ;
        RECT 112.855 64.820 113.385 64.890 ;
        RECT 110.925 64.380 111.925 64.795 ;
        RECT 115.050 64.505 115.220 65.520 ;
        RECT 113.990 64.335 115.220 64.505 ;
        RECT 115.540 64.890 121.120 65.060 ;
        RECT 96.465 63.775 97.060 63.810 ;
        RECT 96.285 63.640 97.060 63.775 ;
        RECT 96.285 63.605 96.815 63.640 ;
        RECT 97.700 63.085 98.700 64.085 ;
        RECT 113.990 63.840 114.160 64.335 ;
        RECT 113.195 62.840 114.195 63.840 ;
        RECT 115.540 63.565 115.710 64.890 ;
        RECT 116.370 64.260 121.120 64.430 ;
        RECT 116.765 63.840 116.935 64.260 ;
        RECT 121.555 64.180 121.885 70.335 ;
        RECT 115.115 63.530 115.710 63.565 ;
        RECT 114.935 63.395 115.710 63.530 ;
        RECT 114.935 63.360 115.465 63.395 ;
        RECT 116.350 62.840 117.350 63.840 ;
        RECT 107.200 57.730 107.865 57.900 ;
        RECT 71.700 55.685 72.000 55.950 ;
        RECT 71.700 55.385 72.245 55.685 ;
        RECT 74.325 55.625 74.855 56.155 ;
        RECT 58.260 54.455 58.790 54.985 ;
        RECT 51.840 54.305 52.010 54.310 ;
        RECT 51.840 54.135 57.620 54.305 ;
        RECT 71.945 54.140 72.245 55.385 ;
        RECT 84.080 54.310 84.380 56.370 ;
        RECT 106.300 56.325 107.300 56.795 ;
        RECT 107.695 56.785 107.865 57.730 ;
        RECT 108.550 57.205 109.550 58.205 ;
        RECT 110.205 57.730 110.985 57.900 ;
        RECT 109.285 56.995 109.455 57.205 ;
        RECT 109.285 56.825 110.490 56.995 ;
        RECT 107.695 56.615 108.955 56.785 ;
        RECT 108.785 56.360 108.955 56.615 ;
        RECT 106.300 56.155 108.440 56.325 ;
        RECT 108.785 56.190 109.995 56.360 ;
        RECT 106.300 55.795 107.300 56.155 ;
        RECT 108.270 55.800 108.440 56.155 ;
        RECT 108.270 55.630 109.470 55.800 ;
        RECT 109.300 55.180 109.470 55.630 ;
        RECT 109.825 55.690 109.995 56.190 ;
        RECT 110.320 56.205 110.490 56.825 ;
        RECT 110.815 56.725 110.985 57.730 ;
        RECT 111.550 57.790 112.550 58.205 ;
        RECT 111.550 57.205 112.620 57.790 ;
        RECT 110.815 56.555 112.150 56.725 ;
        RECT 110.320 56.035 111.670 56.205 ;
        RECT 109.825 55.520 111.210 55.690 ;
        RECT 84.080 54.140 84.410 54.310 ;
        RECT 51.840 53.695 52.010 54.135 ;
        RECT 51.380 52.695 52.380 53.695 ;
        RECT 71.830 53.610 72.360 54.140 ;
        RECT 83.985 53.610 84.515 54.140 ;
        RECT 105.965 54.120 106.965 55.120 ;
        RECT 109.300 55.010 110.695 55.180 ;
        RECT 107.755 54.655 108.820 54.825 ;
        RECT 108.650 54.585 108.820 54.655 ;
        RECT 108.650 54.415 110.195 54.585 ;
        RECT 106.635 53.775 106.805 54.120 ;
        RECT 51.095 51.625 52.185 51.955 ;
        RECT 60.010 51.910 60.900 52.800 ;
        RECT 64.140 52.245 64.870 52.250 ;
        RECT 63.960 52.235 64.870 52.245 ;
        RECT 63.960 52.080 71.560 52.235 ;
        RECT 63.960 52.075 64.490 52.080 ;
        RECT 64.770 52.065 71.560 52.080 ;
        RECT 51.095 47.415 51.425 51.625 ;
        RECT 51.655 51.585 52.185 51.625 ;
        RECT 51.850 50.945 52.020 51.585 ;
        RECT 61.395 51.325 62.395 51.805 ;
        RECT 61.395 51.155 71.560 51.325 ;
        RECT 51.850 50.775 57.620 50.945 ;
        RECT 61.395 50.805 62.395 51.155 ;
        RECT 64.140 50.425 65.000 50.430 ;
        RECT 63.960 50.415 65.000 50.425 ;
        RECT 63.960 50.260 71.560 50.415 ;
        RECT 63.960 50.255 64.490 50.260 ;
        RECT 64.770 50.245 71.560 50.260 ;
        RECT 61.395 49.505 62.395 49.920 ;
        RECT 58.280 48.885 58.810 49.415 ;
        RECT 61.395 49.335 71.560 49.505 ;
        RECT 61.395 48.920 62.395 49.335 ;
        RECT 64.140 48.605 64.980 48.610 ;
        RECT 63.960 48.595 64.980 48.605 ;
        RECT 63.960 48.440 71.560 48.595 ;
        RECT 63.960 48.435 64.490 48.440 ;
        RECT 64.770 48.425 71.560 48.440 ;
        RECT 61.395 47.685 62.395 48.095 ;
        RECT 51.840 47.665 52.010 47.685 ;
        RECT 51.840 47.495 57.620 47.665 ;
        RECT 61.395 47.515 71.560 47.685 ;
        RECT 51.840 47.070 52.010 47.495 ;
        RECT 61.395 47.095 62.395 47.515 ;
        RECT 37.250 45.150 38.500 46.400 ;
        RECT 51.380 46.070 52.380 47.070 ;
        RECT 63.970 46.770 64.500 46.785 ;
        RECT 64.770 46.770 71.560 46.775 ;
        RECT 63.970 46.615 71.560 46.770 ;
        RECT 64.150 46.605 71.560 46.615 ;
        RECT 64.150 46.600 64.870 46.605 ;
        RECT 61.395 45.865 62.395 46.220 ;
        RECT 61.395 45.695 71.560 45.865 ;
        RECT 43.820 45.285 44.350 45.455 ;
        RECT 37.625 44.825 37.925 45.150 ;
        RECT 37.625 41.215 37.955 44.825 ;
        RECT 43.995 44.745 44.165 45.285 ;
        RECT 48.395 45.280 48.925 45.450 ;
        RECT 38.430 44.575 44.200 44.745 ;
        RECT 43.995 44.565 44.165 44.575 ;
        RECT 47.750 43.425 48.080 44.825 ;
        RECT 48.570 44.745 48.740 45.280 ;
        RECT 61.395 45.220 62.395 45.695 ;
        RECT 63.970 44.950 64.500 44.965 ;
        RECT 64.770 44.950 71.560 44.955 ;
        RECT 63.970 44.795 71.560 44.950 ;
        RECT 64.150 44.785 71.560 44.795 ;
        RECT 64.150 44.780 64.920 44.785 ;
        RECT 48.555 44.575 54.325 44.745 ;
        RECT 48.570 44.560 48.740 44.575 ;
        RECT 46.995 43.310 48.080 43.425 ;
        RECT 61.395 44.045 62.395 44.400 ;
        RECT 61.395 43.875 71.560 44.045 ;
        RECT 61.395 43.400 62.395 43.875 ;
        RECT 44.980 42.725 45.510 43.255 ;
        RECT 46.895 43.140 48.080 43.310 ;
        RECT 64.150 43.140 65.015 43.150 ;
        RECT 46.995 43.095 48.080 43.140 ;
        RECT 38.430 41.295 44.200 41.465 ;
        RECT 39.765 40.840 39.935 41.295 ;
        RECT 47.750 41.215 48.080 43.095 ;
        RECT 63.970 43.135 65.015 43.140 ;
        RECT 63.970 42.980 71.560 43.135 ;
        RECT 63.970 42.970 64.500 42.980 ;
        RECT 64.770 42.965 71.560 42.980 ;
        RECT 55.040 42.310 55.570 42.840 ;
        RECT 61.395 42.225 62.395 42.660 ;
        RECT 61.395 42.055 71.560 42.225 ;
        RECT 61.395 41.660 62.395 42.055 ;
        RECT 48.555 41.295 54.325 41.465 ;
        RECT 63.960 41.315 65.005 41.330 ;
        RECT 48.575 40.850 48.745 41.295 ;
        RECT 63.960 41.160 71.560 41.315 ;
        RECT 64.770 41.145 71.560 41.160 ;
        RECT 39.305 39.840 40.305 40.840 ;
        RECT 48.115 39.850 49.115 40.850 ;
        RECT 61.395 40.405 62.395 40.825 ;
        RECT 61.395 40.235 71.560 40.405 ;
        RECT 61.395 39.825 62.395 40.235 ;
        RECT 37.250 38.420 38.500 39.670 ;
        RECT 64.235 39.510 64.430 39.625 ;
        RECT 64.235 39.505 64.965 39.510 ;
        RECT 63.970 39.495 64.965 39.505 ;
        RECT 63.970 39.340 71.560 39.495 ;
        RECT 63.970 39.335 64.500 39.340 ;
        RECT 64.770 39.325 71.560 39.340 ;
        RECT 71.975 39.245 72.305 53.610 ;
        RECT 74.650 51.775 75.260 52.445 ;
        RECT 75.650 51.770 76.180 51.950 ;
        RECT 84.080 51.855 84.410 53.610 ;
        RECT 106.635 53.605 109.600 53.775 ;
        RECT 106.895 52.650 108.750 52.655 ;
        RECT 106.715 52.485 108.750 52.650 ;
        RECT 106.715 52.480 107.245 52.485 ;
        RECT 76.890 51.770 83.680 51.775 ;
        RECT 75.650 51.605 83.680 51.770 ;
        RECT 84.080 51.645 84.425 51.855 ;
        RECT 75.650 51.600 77.070 51.605 ;
        RECT 75.650 51.420 76.180 51.600 ;
        RECT 72.930 50.490 73.930 50.920 ;
        RECT 76.890 50.490 83.680 50.495 ;
        RECT 72.930 50.325 83.680 50.490 ;
        RECT 72.930 50.320 77.065 50.325 ;
        RECT 72.930 49.920 73.930 50.320 ;
        RECT 75.575 49.210 76.105 49.385 ;
        RECT 76.890 49.210 83.680 49.215 ;
        RECT 75.575 49.045 83.680 49.210 ;
        RECT 75.575 49.040 76.960 49.045 ;
        RECT 75.575 48.855 76.105 49.040 ;
        RECT 72.870 47.930 73.870 48.350 ;
        RECT 76.890 47.930 83.680 47.935 ;
        RECT 72.870 47.765 83.680 47.930 ;
        RECT 72.870 47.760 76.960 47.765 ;
        RECT 72.870 47.350 73.870 47.760 ;
        RECT 75.570 46.650 76.100 46.830 ;
        RECT 76.890 46.650 83.680 46.655 ;
        RECT 75.570 46.485 83.680 46.650 ;
        RECT 75.570 46.480 76.960 46.485 ;
        RECT 75.570 46.300 76.100 46.480 ;
        RECT 72.980 45.370 73.980 45.845 ;
        RECT 76.890 45.370 83.680 45.375 ;
        RECT 72.980 45.205 83.680 45.370 ;
        RECT 72.980 45.200 76.960 45.205 ;
        RECT 72.980 44.845 73.980 45.200 ;
        RECT 75.610 44.090 76.140 44.265 ;
        RECT 76.890 44.090 83.680 44.095 ;
        RECT 75.610 43.925 83.680 44.090 ;
        RECT 75.610 43.920 76.960 43.925 ;
        RECT 75.610 43.735 76.140 43.920 ;
        RECT 72.980 42.810 73.980 43.235 ;
        RECT 76.890 42.810 83.680 42.815 ;
        RECT 72.980 42.645 83.680 42.810 ;
        RECT 72.980 42.640 76.960 42.645 ;
        RECT 72.980 42.235 73.980 42.640 ;
        RECT 75.585 41.530 76.115 41.705 ;
        RECT 76.890 41.530 83.680 41.535 ;
        RECT 75.585 41.365 83.680 41.530 ;
        RECT 75.585 41.360 76.960 41.365 ;
        RECT 75.585 41.175 76.115 41.360 ;
        RECT 72.980 40.250 73.980 40.750 ;
        RECT 76.890 40.250 83.680 40.255 ;
        RECT 72.980 40.085 83.680 40.250 ;
        RECT 72.980 40.080 76.960 40.085 ;
        RECT 72.980 39.750 73.980 40.080 ;
        RECT 43.840 38.625 44.370 38.795 ;
        RECT 48.395 38.650 48.925 38.820 ;
        RECT 76.890 38.805 83.680 38.975 ;
        RECT 37.630 38.130 37.950 38.420 ;
        RECT 37.625 34.520 37.955 38.130 ;
        RECT 44.015 38.050 44.185 38.625 ;
        RECT 38.430 37.880 44.200 38.050 ;
        RECT 44.950 36.020 45.480 36.550 ;
        RECT 47.750 36.380 48.080 38.130 ;
        RECT 48.570 38.050 48.740 38.650 ;
        RECT 76.060 38.100 76.590 38.280 ;
        RECT 77.650 38.100 77.820 38.805 ;
        RECT 84.095 38.725 84.425 51.645 ;
        RECT 108.580 51.700 108.750 52.485 ;
        RECT 109.430 52.330 109.600 53.605 ;
        RECT 110.025 52.960 110.195 54.415 ;
        RECT 110.525 53.590 110.695 55.010 ;
        RECT 111.040 54.220 111.210 55.520 ;
        RECT 111.500 54.850 111.670 56.035 ;
        RECT 111.980 55.480 112.150 56.555 ;
        RECT 112.450 56.110 112.620 57.205 ;
        RECT 114.090 56.740 114.790 57.900 ;
        RECT 113.535 56.570 120.325 56.740 ;
        RECT 112.450 55.940 120.325 56.110 ;
        RECT 111.980 55.310 120.325 55.480 ;
        RECT 111.500 54.680 120.325 54.850 ;
        RECT 111.040 54.050 120.325 54.220 ;
        RECT 110.525 53.420 120.325 53.590 ;
        RECT 110.025 52.790 120.325 52.960 ;
        RECT 109.430 52.160 120.325 52.330 ;
        RECT 120.740 51.705 121.070 56.820 ;
        RECT 108.580 51.530 120.325 51.700 ;
        RECT 105.965 51.070 106.965 51.500 ;
        RECT 105.965 50.900 120.325 51.070 ;
        RECT 120.740 51.005 122.445 51.705 ;
        RECT 105.965 50.500 106.965 50.900 ;
        RECT 108.420 50.270 120.325 50.440 ;
        RECT 108.420 49.375 108.590 50.270 ;
        RECT 106.895 49.370 108.590 49.375 ;
        RECT 106.715 49.205 108.590 49.370 ;
        RECT 109.310 49.810 113.700 49.820 ;
        RECT 109.310 49.650 120.325 49.810 ;
        RECT 106.715 49.200 107.245 49.205 ;
        RECT 109.310 48.510 109.480 49.650 ;
        RECT 113.535 49.640 120.325 49.650 ;
        RECT 108.515 48.340 109.480 48.510 ;
        RECT 109.920 49.010 120.325 49.180 ;
        RECT 108.515 48.255 108.685 48.340 ;
        RECT 106.380 48.085 108.685 48.255 ;
        RECT 106.380 47.750 106.550 48.085 ;
        RECT 109.920 47.835 110.090 49.010 ;
        RECT 105.965 46.750 106.965 47.750 ;
        RECT 109.125 47.665 110.090 47.835 ;
        RECT 110.445 48.380 120.325 48.550 ;
        RECT 109.125 47.330 109.295 47.665 ;
        RECT 107.755 47.160 109.295 47.330 ;
        RECT 110.445 47.215 110.615 48.380 ;
        RECT 109.665 47.045 110.615 47.215 ;
        RECT 111.030 47.750 120.325 47.920 ;
        RECT 109.665 46.215 109.835 47.045 ;
        RECT 111.030 46.635 111.200 47.750 ;
        RECT 106.640 45.660 107.640 46.145 ;
        RECT 108.675 46.045 109.835 46.215 ;
        RECT 110.205 46.465 111.200 46.635 ;
        RECT 111.520 47.120 120.325 47.290 ;
        RECT 108.675 45.660 108.845 46.045 ;
        RECT 106.640 45.490 108.845 45.660 ;
        RECT 110.205 45.635 110.375 46.465 ;
        RECT 111.520 46.025 111.690 47.120 ;
        RECT 106.640 45.145 107.640 45.490 ;
        RECT 109.340 45.465 110.375 45.635 ;
        RECT 110.725 45.855 111.690 46.025 ;
        RECT 112.080 46.490 120.325 46.660 ;
        RECT 109.340 45.200 109.510 45.465 ;
        RECT 108.250 45.030 109.510 45.200 ;
        RECT 110.725 45.150 110.895 45.855 ;
        RECT 112.080 45.385 112.250 46.490 ;
        RECT 108.250 44.200 108.420 45.030 ;
        RECT 109.890 44.980 110.895 45.150 ;
        RECT 111.235 45.215 112.250 45.385 ;
        RECT 112.740 45.860 120.325 46.030 ;
        RECT 109.890 44.655 110.060 44.980 ;
        RECT 107.755 44.030 108.420 44.200 ;
        RECT 107.935 44.020 108.420 44.030 ;
        RECT 109.050 44.070 110.060 44.655 ;
        RECT 111.235 44.200 111.405 45.215 ;
        RECT 112.740 44.695 112.910 45.860 ;
        RECT 113.535 45.230 120.325 45.400 ;
        RECT 114.345 45.225 114.525 45.230 ;
        RECT 110.835 44.175 111.405 44.200 ;
        RECT 109.050 43.655 110.050 44.070 ;
        RECT 110.655 44.030 111.405 44.175 ;
        RECT 111.780 44.125 112.910 44.695 ;
        RECT 114.355 44.430 114.525 45.225 ;
        RECT 120.740 45.150 121.070 51.005 ;
        RECT 114.175 44.260 114.705 44.430 ;
        RECT 110.655 44.005 111.185 44.030 ;
        RECT 111.780 43.695 112.780 44.125 ;
        RECT 112.765 41.665 113.295 42.195 ;
        RECT 48.555 37.880 54.325 38.050 ;
        RECT 76.060 37.930 77.820 38.100 ;
        RECT 76.060 37.750 76.590 37.930 ;
        RECT 57.855 36.505 58.385 36.835 ;
        RECT 46.995 36.345 48.080 36.380 ;
        RECT 46.895 36.175 48.080 36.345 ;
        RECT 46.995 36.050 48.080 36.175 ;
        RECT 38.430 34.600 44.200 34.770 ;
        RECT 39.415 34.135 39.585 34.600 ;
        RECT 47.750 34.520 48.080 36.050 ;
        RECT 55.060 35.975 55.590 36.505 ;
        RECT 58.055 35.150 58.385 36.505 ;
        RECT 58.955 35.615 59.955 36.615 ;
        RECT 72.850 36.030 73.740 36.920 ;
        RECT 58.655 35.150 58.985 35.195 ;
        RECT 58.055 34.820 58.985 35.150 ;
        RECT 59.455 35.115 59.625 35.615 ;
        RECT 59.400 34.945 66.190 35.115 ;
        RECT 48.555 34.600 54.325 34.770 ;
        RECT 48.560 34.145 48.730 34.600 ;
        RECT 37.250 32.325 38.500 33.575 ;
        RECT 38.955 33.135 39.955 34.135 ;
        RECT 48.100 33.145 49.100 34.145 ;
        RECT 58.655 33.955 58.985 34.820 ;
        RECT 66.560 34.255 67.170 34.925 ;
        RECT 72.105 34.900 72.435 35.370 ;
        RECT 73.285 35.290 73.455 36.030 ;
        RECT 72.850 35.120 79.640 35.290 ;
        RECT 71.035 34.840 72.435 34.900 ;
        RECT 70.935 34.670 72.435 34.840 ;
        RECT 71.035 34.570 72.435 34.670 ;
        RECT 59.400 34.035 66.190 34.205 ;
        RECT 72.105 34.130 72.435 34.570 ;
        RECT 72.850 34.210 79.640 34.380 ;
        RECT 80.610 34.375 81.220 35.045 ;
        RECT 59.415 33.570 59.585 34.035 ;
        RECT 43.800 32.510 44.330 32.680 ;
        RECT 37.635 32.015 37.955 32.325 ;
        RECT 37.625 28.405 37.955 32.015 ;
        RECT 43.975 31.935 44.145 32.510 ;
        RECT 49.585 32.490 50.115 32.660 ;
        RECT 58.955 32.570 59.955 33.570 ;
        RECT 73.495 33.490 73.665 34.210 ;
        RECT 73.315 32.960 73.845 33.490 ;
        RECT 38.430 31.765 44.200 31.935 ;
        RECT 44.950 29.930 45.480 30.460 ;
        RECT 47.750 30.140 48.080 32.015 ;
        RECT 49.760 31.935 49.930 32.490 ;
        RECT 48.555 31.765 54.325 31.935 ;
        RECT 46.895 29.810 48.080 30.140 ;
        RECT 55.060 29.950 55.590 30.480 ;
        RECT 38.430 28.485 44.200 28.655 ;
        RECT 39.415 28.020 39.585 28.485 ;
        RECT 47.750 28.405 48.080 29.810 ;
        RECT 48.595 28.655 48.765 28.665 ;
        RECT 48.555 28.485 54.325 28.655 ;
        RECT 48.595 28.050 48.765 28.485 ;
        RECT 37.420 25.955 38.670 27.205 ;
        RECT 38.955 27.020 39.955 28.020 ;
        RECT 48.135 27.050 49.135 28.050 ;
        RECT 63.515 27.570 63.685 28.240 ;
        RECT 43.840 26.085 44.370 26.255 ;
        RECT 49.585 26.085 50.115 26.255 ;
        RECT 37.640 25.610 37.940 25.955 ;
        RECT 37.625 22.000 37.955 25.610 ;
        RECT 44.015 25.530 44.185 26.085 ;
        RECT 38.430 25.360 44.200 25.530 ;
        RECT 47.750 24.055 48.080 25.610 ;
        RECT 49.760 25.530 49.930 26.085 ;
        RECT 48.555 25.360 54.325 25.530 ;
        RECT 63.515 25.150 63.685 27.030 ;
        RECT 88.580 26.360 88.750 28.240 ;
        RECT 46.995 23.985 48.080 24.055 ;
        RECT 44.950 23.455 45.480 23.985 ;
        RECT 46.895 23.815 48.080 23.985 ;
        RECT 46.995 23.725 48.080 23.815 ;
        RECT 38.430 22.240 44.200 22.250 ;
        RECT 38.425 22.080 44.200 22.240 ;
        RECT 38.425 21.625 38.595 22.080 ;
        RECT 47.750 22.000 48.080 23.725 ;
        RECT 55.060 23.605 55.590 24.135 ;
        RECT 63.515 22.730 63.685 24.610 ;
        RECT 88.580 23.940 88.750 25.820 ;
        RECT 88.580 22.730 88.750 23.400 ;
        RECT 48.550 22.250 48.720 22.260 ;
        RECT 48.550 22.080 54.325 22.250 ;
        RECT 48.550 21.645 48.720 22.080 ;
        RECT 37.965 20.625 38.965 21.625 ;
        RECT 48.090 20.645 49.090 21.645 ;
      LAYER mcon ;
        RECT 53.695 209.790 54.225 210.320 ;
        RECT 97.395 210.305 97.565 210.475 ;
        RECT 97.755 210.305 97.925 210.475 ;
        RECT 51.665 207.770 52.195 208.300 ;
        RECT 105.590 210.445 105.760 210.615 ;
        RECT 105.950 210.445 106.120 210.615 ;
        RECT 53.685 204.725 54.215 205.255 ;
        RECT 51.665 202.870 52.195 203.400 ;
        RECT 97.395 203.130 97.565 203.300 ;
        RECT 97.755 203.130 97.925 203.300 ;
        RECT 105.590 203.365 105.760 203.535 ;
        RECT 105.950 203.365 106.120 203.535 ;
        RECT 81.320 199.665 81.850 200.195 ;
        RECT 53.610 198.295 54.140 198.825 ;
        RECT 83.145 198.335 83.675 198.865 ;
        RECT 51.665 196.335 52.195 196.865 ;
        RECT 104.385 197.270 104.915 197.800 ;
        RECT 112.465 197.270 112.995 197.800 ;
        RECT 97.395 196.180 97.565 196.350 ;
        RECT 97.755 196.180 97.925 196.350 ;
        RECT 53.665 193.370 54.195 193.900 ;
        RECT 105.590 196.495 105.760 196.665 ;
        RECT 105.950 196.495 106.120 196.665 ;
        RECT 51.665 191.645 52.195 192.175 ;
        RECT 81.320 192.560 81.850 193.090 ;
        RECT 83.145 191.435 83.675 191.965 ;
        RECT 104.385 190.205 104.915 190.735 ;
        RECT 97.395 189.155 97.565 189.325 ;
        RECT 97.755 189.155 97.925 189.325 ;
        RECT 112.465 189.765 112.995 190.295 ;
        RECT 105.590 189.155 105.760 189.325 ;
        RECT 105.950 189.155 106.120 189.325 ;
        RECT 46.430 185.335 46.960 185.865 ;
        RECT 44.420 184.075 44.950 184.605 ;
        RECT 58.315 182.800 58.485 182.970 ;
        RECT 58.315 182.440 58.485 182.610 ;
        RECT 118.650 182.800 118.820 182.970 ;
        RECT 118.650 182.440 118.820 182.610 ;
        RECT 58.315 181.590 58.485 181.760 ;
        RECT 58.315 181.230 58.485 181.400 ;
        RECT 118.650 181.590 118.820 181.760 ;
        RECT 118.650 181.230 118.820 181.400 ;
        RECT 46.430 180.605 46.960 181.135 ;
        RECT 58.315 180.380 58.485 180.550 ;
        RECT 44.420 179.620 44.950 180.150 ;
        RECT 58.315 180.020 58.485 180.190 ;
        RECT 118.650 180.380 118.820 180.550 ;
        RECT 118.650 180.020 118.820 180.190 ;
        RECT 58.315 179.170 58.485 179.340 ;
        RECT 58.315 178.810 58.485 178.980 ;
        RECT 118.650 179.170 118.820 179.340 ;
        RECT 118.650 178.810 118.820 178.980 ;
        RECT 58.315 177.960 58.485 178.130 ;
        RECT 58.315 177.600 58.485 177.770 ;
        RECT 118.650 177.960 118.820 178.130 ;
        RECT 118.650 177.600 118.820 177.770 ;
        RECT 58.315 176.750 58.485 176.920 ;
        RECT 46.430 176.040 46.960 176.570 ;
        RECT 58.315 176.390 58.485 176.560 ;
        RECT 118.650 176.750 118.820 176.920 ;
        RECT 118.650 176.390 118.820 176.560 ;
        RECT 44.420 175.020 44.950 175.550 ;
        RECT 106.855 173.225 107.385 173.755 ;
        RECT 46.345 170.470 46.875 171.000 ;
        RECT 112.970 171.460 113.500 171.990 ;
        RECT 90.960 170.795 91.490 171.325 ;
        RECT 44.420 169.475 44.950 170.005 ;
        RECT 105.560 170.090 105.730 170.260 ;
        RECT 105.920 170.090 106.090 170.260 ;
        RECT 107.075 167.400 107.605 167.930 ;
        RECT 52.385 166.635 52.915 167.165 ;
        RECT 46.345 166.020 46.875 166.550 ;
        RECT 106.855 166.055 107.385 166.585 ;
        RECT 44.485 164.835 45.015 165.365 ;
        RECT 112.880 164.905 113.410 165.435 ;
        RECT 105.560 163.300 105.730 163.470 ;
        RECT 105.920 163.300 106.090 163.470 ;
        RECT 52.320 162.000 52.850 162.530 ;
        RECT 46.345 161.445 46.875 161.975 ;
        RECT 44.420 160.370 44.950 160.900 ;
        RECT 91.025 160.865 91.555 161.395 ;
        RECT 107.075 160.270 107.605 160.800 ;
        RECT 52.325 157.250 52.855 157.780 ;
        RECT 45.675 155.140 45.845 155.310 ;
        RECT 45.675 154.780 45.845 154.950 ;
        RECT 110.680 155.140 110.850 155.310 ;
        RECT 110.680 154.780 110.850 154.950 ;
        RECT 45.675 153.930 45.845 154.100 ;
        RECT 45.675 153.570 45.845 153.740 ;
        RECT 110.680 153.930 110.850 154.100 ;
        RECT 110.680 153.570 110.850 153.740 ;
        RECT 45.675 152.720 45.845 152.890 ;
        RECT 45.675 152.360 45.845 152.530 ;
        RECT 110.680 152.720 110.850 152.890 ;
        RECT 110.680 152.360 110.850 152.530 ;
        RECT 45.675 151.510 45.845 151.680 ;
        RECT 45.675 151.150 45.845 151.320 ;
        RECT 110.680 151.510 110.850 151.680 ;
        RECT 110.680 151.150 110.850 151.320 ;
        RECT 45.675 150.300 45.845 150.470 ;
        RECT 45.675 149.940 45.845 150.110 ;
        RECT 110.680 150.300 110.850 150.470 ;
        RECT 110.680 149.940 110.850 150.110 ;
        RECT 45.675 149.090 45.845 149.260 ;
        RECT 45.675 148.730 45.845 148.900 ;
        RECT 110.680 149.090 110.850 149.260 ;
        RECT 110.680 148.730 110.850 148.900 ;
        RECT 45.675 147.880 45.845 148.050 ;
        RECT 45.675 147.520 45.845 147.690 ;
        RECT 110.680 147.880 110.850 148.050 ;
        RECT 110.680 147.520 110.850 147.690 ;
        RECT 45.675 146.670 45.845 146.840 ;
        RECT 45.675 146.310 45.845 146.480 ;
        RECT 110.680 146.670 110.850 146.840 ;
        RECT 110.680 146.310 110.850 146.480 ;
        RECT 45.675 145.460 45.845 145.630 ;
        RECT 45.675 145.100 45.845 145.270 ;
        RECT 110.680 145.460 110.850 145.630 ;
        RECT 110.680 145.100 110.850 145.270 ;
        RECT 45.675 144.250 45.845 144.420 ;
        RECT 45.675 143.890 45.845 144.060 ;
        RECT 110.680 144.250 110.850 144.420 ;
        RECT 110.680 143.890 110.850 144.060 ;
        RECT 45.675 143.040 45.845 143.210 ;
        RECT 45.675 142.680 45.845 142.850 ;
        RECT 110.680 143.040 110.850 143.210 ;
        RECT 110.680 142.680 110.850 142.850 ;
        RECT 45.675 141.830 45.845 142.000 ;
        RECT 45.675 141.470 45.845 141.640 ;
        RECT 110.680 141.830 110.850 142.000 ;
        RECT 110.680 141.470 110.850 141.640 ;
        RECT 45.675 140.620 45.845 140.790 ;
        RECT 45.675 140.260 45.845 140.430 ;
        RECT 110.680 140.620 110.850 140.790 ;
        RECT 110.680 140.260 110.850 140.430 ;
        RECT 45.675 139.410 45.845 139.580 ;
        RECT 45.675 139.050 45.845 139.220 ;
        RECT 110.680 139.410 110.850 139.580 ;
        RECT 110.680 139.050 110.850 139.220 ;
        RECT 45.675 138.200 45.845 138.370 ;
        RECT 45.675 137.840 45.845 138.010 ;
        RECT 110.680 138.200 110.850 138.370 ;
        RECT 110.680 137.840 110.850 138.010 ;
        RECT 45.675 136.990 45.845 137.160 ;
        RECT 45.675 136.630 45.845 136.800 ;
        RECT 110.680 136.990 110.850 137.160 ;
        RECT 110.680 136.630 110.850 136.800 ;
        RECT 78.770 109.435 78.940 109.605 ;
        RECT 79.130 109.435 79.300 109.605 ;
        RECT 46.405 108.900 46.575 109.070 ;
        RECT 55.390 108.910 55.560 109.080 ;
        RECT 65.625 108.910 65.795 109.080 ;
        RECT 44.290 106.385 44.460 106.555 ;
        RECT 44.650 106.385 44.820 106.555 ;
        RECT 61.505 106.240 61.675 106.410 ;
        RECT 61.865 106.240 62.035 106.410 ;
        RECT 71.530 106.240 71.700 106.410 ;
        RECT 71.890 106.240 72.060 106.410 ;
        RECT 45.840 102.555 46.730 103.085 ;
        RECT 54.825 102.590 55.715 103.120 ;
        RECT 65.320 102.530 66.210 103.060 ;
        RECT 82.960 104.845 83.130 105.015 ;
        RECT 82.960 104.485 83.130 104.655 ;
        RECT 123.795 104.845 123.965 105.015 ;
        RECT 123.795 104.485 123.965 104.655 ;
        RECT 79.780 102.525 79.950 102.695 ;
        RECT 82.960 103.635 83.130 103.805 ;
        RECT 82.960 103.275 83.130 103.445 ;
        RECT 123.795 103.635 123.965 103.805 ;
        RECT 123.795 103.275 123.965 103.445 ;
        RECT 82.960 102.425 83.130 102.595 ;
        RECT 82.960 102.065 83.130 102.235 ;
        RECT 123.795 102.425 123.965 102.595 ;
        RECT 123.795 102.065 123.965 102.235 ;
        RECT 82.960 101.215 83.130 101.385 ;
        RECT 82.960 100.855 83.130 101.025 ;
        RECT 46.405 100.050 46.575 100.220 ;
        RECT 123.795 101.215 123.965 101.385 ;
        RECT 123.795 100.855 123.965 101.025 ;
        RECT 82.960 100.005 83.130 100.175 ;
        RECT 78.695 99.435 78.865 99.605 ;
        RECT 79.055 99.435 79.225 99.605 ;
        RECT 82.960 99.645 83.130 99.815 ;
        RECT 123.795 100.005 123.965 100.175 ;
        RECT 123.795 99.645 123.965 99.815 ;
        RECT 55.390 98.950 55.560 99.120 ;
        RECT 65.625 98.970 65.795 99.140 ;
        RECT 44.290 96.590 44.460 96.760 ;
        RECT 44.650 96.590 44.820 96.760 ;
        RECT 61.505 95.890 61.675 96.060 ;
        RECT 61.865 95.890 62.035 96.060 ;
        RECT 71.530 95.890 71.700 96.060 ;
        RECT 71.890 95.890 72.060 96.060 ;
        RECT 45.840 92.645 46.730 93.175 ;
        RECT 54.825 92.680 55.715 93.210 ;
        RECT 65.320 92.635 66.210 93.165 ;
        RECT 96.510 95.855 97.400 96.385 ;
        RECT 98.505 95.840 98.675 96.010 ;
        RECT 114.840 95.855 115.730 96.385 ;
        RECT 94.605 94.130 95.495 94.660 ;
        RECT 96.575 94.590 96.745 94.760 ;
        RECT 79.780 93.005 79.950 93.175 ;
        RECT 93.575 92.565 94.465 93.095 ;
        RECT 116.835 95.840 117.005 96.010 ;
        RECT 104.640 93.445 105.530 93.975 ;
        RECT 112.935 94.130 113.825 94.660 ;
        RECT 114.905 94.590 115.075 94.760 ;
        RECT 95.525 92.920 95.695 93.090 ;
        RECT 91.225 91.060 92.115 91.590 ;
        RECT 93.410 91.340 93.580 91.510 ;
        RECT 89.850 90.525 90.020 90.695 ;
        RECT 90.210 90.525 90.380 90.695 ;
        RECT 78.695 89.605 78.865 89.775 ;
        RECT 79.055 89.605 79.225 89.775 ;
        RECT 55.390 89.180 55.560 89.350 ;
        RECT 65.625 89.305 65.795 89.475 ;
        RECT 46.405 88.830 46.575 89.000 ;
        RECT 44.290 87.230 44.460 87.400 ;
        RECT 44.650 87.230 44.820 87.400 ;
        RECT 88.010 88.900 88.900 89.430 ;
        RECT 61.505 85.870 61.675 86.040 ;
        RECT 61.865 85.870 62.035 86.040 ;
        RECT 71.530 86.030 71.700 86.200 ;
        RECT 71.890 86.030 72.060 86.200 ;
        RECT 45.840 82.490 46.730 83.020 ;
        RECT 54.825 82.665 55.715 83.195 ;
        RECT 65.320 82.780 66.210 83.310 ;
        RECT 74.365 82.930 75.255 83.460 ;
        RECT 90.210 88.165 90.380 88.335 ;
        RECT 90.545 86.520 91.435 87.050 ;
        RECT 92.545 86.700 92.715 86.870 ;
        RECT 92.620 85.095 93.510 85.625 ;
        RECT 94.650 85.180 94.820 85.350 ;
        RECT 92.620 83.150 93.510 83.680 ;
        RECT 94.855 83.355 95.025 83.525 ;
        RECT 79.745 82.650 79.915 82.820 ;
        RECT 94.890 81.610 95.780 82.140 ;
        RECT 111.905 92.565 112.795 93.095 ;
        RECT 113.855 92.920 114.025 93.090 ;
        RECT 109.555 91.060 110.445 91.590 ;
        RECT 111.740 91.340 111.910 91.510 ;
        RECT 108.180 90.525 108.350 90.695 ;
        RECT 108.540 90.525 108.710 90.695 ;
        RECT 106.340 88.920 107.230 89.450 ;
        RECT 122.465 89.025 122.995 89.555 ;
        RECT 108.540 88.165 108.710 88.335 ;
        RECT 108.875 86.520 109.765 87.050 ;
        RECT 110.875 86.700 111.045 86.870 ;
        RECT 110.950 85.095 111.840 85.625 ;
        RECT 112.980 85.180 113.150 85.350 ;
        RECT 110.950 83.150 111.840 83.680 ;
        RECT 113.185 83.355 113.355 83.525 ;
        RECT 96.935 81.895 97.105 82.065 ;
        RECT 98.045 81.610 98.935 82.140 ;
        RECT 113.220 81.610 114.110 82.140 ;
        RECT 115.265 81.895 115.435 82.065 ;
        RECT 116.375 81.610 117.265 82.140 ;
        RECT 46.405 79.755 46.575 79.925 ;
        RECT 55.390 79.745 55.560 79.915 ;
        RECT 65.625 79.790 65.795 79.960 ;
        RECT 78.855 79.480 79.025 79.650 ;
        RECT 79.215 79.480 79.385 79.650 ;
        RECT 43.685 76.745 43.855 76.915 ;
        RECT 44.045 76.745 44.215 76.915 ;
        RECT 61.505 76.935 61.675 77.105 ;
        RECT 61.865 76.935 62.035 77.105 ;
        RECT 71.530 76.705 71.700 76.875 ;
        RECT 71.890 76.705 72.060 76.875 ;
        RECT 45.840 73.485 46.730 74.015 ;
        RECT 54.825 73.460 55.715 73.990 ;
        RECT 65.320 73.605 66.210 74.135 ;
        RECT 73.960 73.305 74.850 73.835 ;
        RECT 96.270 77.565 97.160 78.095 ;
        RECT 98.215 77.550 98.385 77.720 ;
        RECT 94.315 75.840 95.205 76.370 ;
        RECT 96.285 76.300 96.455 76.470 ;
        RECT 93.285 74.275 94.175 74.805 ;
        RECT 114.870 77.320 115.760 77.850 ;
        RECT 116.865 77.305 117.035 77.475 ;
        RECT 95.235 74.630 95.405 74.800 ;
        RECT 79.515 73.130 79.685 73.300 ;
        RECT 79.875 73.130 80.045 73.300 ;
        RECT 90.935 72.770 91.825 73.300 ;
        RECT 93.120 73.050 93.290 73.220 ;
        RECT 89.560 72.235 89.730 72.405 ;
        RECT 89.920 72.235 90.090 72.405 ;
        RECT 51.730 71.750 51.900 71.920 ;
        RECT 52.090 71.750 52.260 71.920 ;
        RECT 87.720 70.630 88.610 71.160 ;
        RECT 89.920 69.875 90.090 70.045 ;
        RECT 64.085 68.780 64.255 68.950 ;
        RECT 51.435 66.285 52.325 66.815 ;
        RECT 64.085 66.960 64.255 67.130 ;
        RECT 51.730 65.210 51.900 65.380 ;
        RECT 52.090 65.210 52.260 65.380 ;
        RECT 64.085 65.140 64.255 65.310 ;
        RECT 64.095 63.325 64.265 63.495 ;
        RECT 64.095 61.500 64.265 61.670 ;
        RECT 51.435 59.595 52.325 60.125 ;
        RECT 64.095 59.675 64.265 59.845 ;
        RECT 51.730 58.515 51.900 58.685 ;
        RECT 52.090 58.515 52.260 58.685 ;
        RECT 64.085 57.865 64.255 58.035 ;
        RECT 61.790 56.040 61.960 56.210 ;
        RECT 64.095 56.040 64.265 56.210 ;
        RECT 90.255 68.230 91.145 68.760 ;
        RECT 92.255 68.410 92.425 68.580 ;
        RECT 92.330 66.805 93.220 67.335 ;
        RECT 94.360 66.890 94.530 67.060 ;
        RECT 92.330 64.860 93.220 65.390 ;
        RECT 94.565 65.065 94.735 65.235 ;
        RECT 112.965 75.595 113.855 76.125 ;
        RECT 114.935 76.055 115.105 76.225 ;
        RECT 111.935 74.030 112.825 74.560 ;
        RECT 113.885 74.385 114.055 74.555 ;
        RECT 109.585 72.525 110.475 73.055 ;
        RECT 111.770 72.805 111.940 72.975 ;
        RECT 108.210 71.990 108.380 72.160 ;
        RECT 108.570 71.990 108.740 72.160 ;
        RECT 106.370 70.400 107.260 70.930 ;
        RECT 122.190 70.420 122.720 70.950 ;
        RECT 108.570 69.630 108.740 69.800 ;
        RECT 108.905 67.985 109.795 68.515 ;
        RECT 110.905 68.165 111.075 68.335 ;
        RECT 110.980 66.560 111.870 67.090 ;
        RECT 113.010 66.645 113.180 66.815 ;
        RECT 94.600 63.320 95.490 63.850 ;
        RECT 110.980 64.615 111.870 65.145 ;
        RECT 113.215 64.820 113.385 64.990 ;
        RECT 96.645 63.605 96.815 63.775 ;
        RECT 97.755 63.320 98.645 63.850 ;
        RECT 113.250 63.075 114.140 63.605 ;
        RECT 115.295 63.360 115.465 63.530 ;
        RECT 116.405 63.075 117.295 63.605 ;
        RECT 107.560 57.730 107.730 57.900 ;
        RECT 108.605 57.440 109.495 57.970 ;
        RECT 110.565 57.730 110.735 57.900 ;
        RECT 106.355 56.030 107.245 56.560 ;
        RECT 111.605 57.440 112.495 57.970 ;
        RECT 106.020 54.355 106.910 54.885 ;
        RECT 108.115 54.655 108.285 54.825 ;
        RECT 51.435 52.930 52.325 53.460 ;
        RECT 64.320 52.075 64.490 52.245 ;
        RECT 52.015 51.585 52.185 51.755 ;
        RECT 61.450 51.040 62.340 51.570 ;
        RECT 64.320 50.255 64.490 50.425 ;
        RECT 61.450 49.155 62.340 49.685 ;
        RECT 64.320 48.435 64.490 48.605 ;
        RECT 61.450 47.330 62.340 47.860 ;
        RECT 51.435 46.305 52.325 46.835 ;
        RECT 64.330 46.615 64.500 46.785 ;
        RECT 61.450 45.455 62.340 45.985 ;
        RECT 44.180 45.285 44.350 45.455 ;
        RECT 48.755 45.280 48.925 45.450 ;
        RECT 64.330 44.795 64.500 44.965 ;
        RECT 61.450 43.635 62.340 44.165 ;
        RECT 47.255 43.140 47.425 43.310 ;
        RECT 64.330 42.970 64.500 43.140 ;
        RECT 61.450 41.895 62.340 42.425 ;
        RECT 64.320 41.160 64.490 41.330 ;
        RECT 39.360 40.075 40.250 40.605 ;
        RECT 48.170 40.085 49.060 40.615 ;
        RECT 61.450 40.060 62.340 40.590 ;
        RECT 64.330 39.335 64.500 39.505 ;
        RECT 74.690 51.845 75.220 52.375 ;
        RECT 107.075 52.480 107.245 52.650 ;
        RECT 72.985 50.155 73.875 50.685 ;
        RECT 72.925 47.585 73.815 48.115 ;
        RECT 73.035 45.080 73.925 45.610 ;
        RECT 73.035 42.470 73.925 43.000 ;
        RECT 73.035 39.985 73.925 40.515 ;
        RECT 44.200 38.625 44.370 38.795 ;
        RECT 48.755 38.650 48.925 38.820 ;
        RECT 114.175 57.730 114.345 57.900 ;
        RECT 114.535 57.730 114.705 57.900 ;
        RECT 106.020 50.735 106.910 51.265 ;
        RECT 121.830 51.130 122.360 51.660 ;
        RECT 107.075 49.200 107.245 49.370 ;
        RECT 106.020 46.985 106.910 47.515 ;
        RECT 108.115 47.160 108.285 47.330 ;
        RECT 106.695 45.380 107.585 45.910 ;
        RECT 108.115 44.030 108.285 44.200 ;
        RECT 109.105 43.890 109.995 44.420 ;
        RECT 111.015 44.005 111.185 44.175 ;
        RECT 111.835 43.930 112.725 44.460 ;
        RECT 114.535 44.260 114.705 44.430 ;
        RECT 57.855 36.585 58.025 36.755 ;
        RECT 58.215 36.585 58.385 36.755 ;
        RECT 47.255 36.175 47.425 36.345 ;
        RECT 59.010 35.850 59.900 36.380 ;
        RECT 39.010 33.370 39.900 33.900 ;
        RECT 66.600 34.325 67.130 34.855 ;
        RECT 71.295 34.670 71.465 34.840 ;
        RECT 80.650 34.445 81.180 34.975 ;
        RECT 48.155 33.380 49.045 33.910 ;
        RECT 59.010 32.805 59.900 33.335 ;
        RECT 44.160 32.510 44.330 32.680 ;
        RECT 49.945 32.490 50.115 32.660 ;
        RECT 46.895 29.890 47.065 30.060 ;
        RECT 47.255 29.890 47.425 30.060 ;
        RECT 39.010 27.255 39.900 27.785 ;
        RECT 48.190 27.285 49.080 27.815 ;
        RECT 63.515 28.000 63.685 28.170 ;
        RECT 63.515 27.640 63.685 27.810 ;
        RECT 88.580 28.000 88.750 28.170 ;
        RECT 88.580 27.640 88.750 27.810 ;
        RECT 63.515 26.790 63.685 26.960 ;
        RECT 63.515 26.430 63.685 26.600 ;
        RECT 44.200 26.085 44.370 26.255 ;
        RECT 49.945 26.085 50.115 26.255 ;
        RECT 88.580 26.790 88.750 26.960 ;
        RECT 88.580 26.430 88.750 26.600 ;
        RECT 63.515 25.580 63.685 25.750 ;
        RECT 63.515 25.220 63.685 25.390 ;
        RECT 88.580 25.580 88.750 25.750 ;
        RECT 88.580 25.220 88.750 25.390 ;
        RECT 63.515 24.370 63.685 24.540 ;
        RECT 47.255 23.815 47.425 23.985 ;
        RECT 63.515 24.010 63.685 24.180 ;
        RECT 88.580 24.370 88.750 24.540 ;
        RECT 88.580 24.010 88.750 24.180 ;
        RECT 63.515 23.160 63.685 23.330 ;
        RECT 63.515 22.800 63.685 22.970 ;
        RECT 88.580 23.160 88.750 23.330 ;
        RECT 88.580 22.800 88.750 22.970 ;
        RECT 38.020 20.860 38.910 21.390 ;
        RECT 48.145 20.880 49.035 21.410 ;
      LAYER met1 ;
        RECT 59.870 219.520 88.935 219.590 ;
        RECT 59.825 218.620 88.935 219.520 ;
        RECT 59.870 218.590 88.935 218.620 ;
        RECT 59.870 216.045 60.870 218.590 ;
        RECT 87.935 216.045 88.935 218.590 ;
        RECT 37.425 214.655 43.100 216.045 ;
        RECT 10.685 213.655 43.100 214.655 ;
        RECT 37.425 210.405 43.100 213.655 ;
        RECT 56.045 210.545 66.045 216.045 ;
        RECT 83.785 210.635 93.785 216.045 ;
        RECT 119.920 215.935 124.425 216.045 ;
        RECT 119.920 214.935 128.510 215.935 ;
        RECT 95.500 213.755 114.430 214.455 ;
        RECT 37.425 209.705 54.255 210.405 ;
        RECT 37.425 185.950 43.100 209.705 ;
        RECT 51.470 208.385 52.170 209.705 ;
        RECT 51.470 207.685 52.225 208.385 ;
        RECT 51.490 205.340 52.190 207.685 ;
        RECT 58.740 207.480 59.330 208.130 ;
        RECT 53.265 205.760 53.855 206.410 ;
        RECT 51.490 204.640 54.245 205.340 ;
        RECT 51.490 203.485 52.190 204.640 ;
        RECT 51.490 202.785 52.225 203.485 ;
        RECT 58.885 203.475 59.185 207.480 ;
        RECT 62.425 205.990 63.125 210.545 ;
        RECT 63.840 206.690 64.430 207.340 ;
        RECT 91.335 205.990 92.035 210.635 ;
        RECT 92.925 206.690 93.515 207.340 ;
        RECT 62.300 204.980 63.250 205.990 ;
        RECT 91.210 204.980 92.160 205.990 ;
        RECT 58.740 202.825 59.330 203.475 ;
        RECT 63.660 202.885 64.250 203.535 ;
        RECT 92.925 202.905 93.515 203.555 ;
        RECT 51.510 198.910 52.210 202.785 ;
        RECT 53.225 200.950 53.815 201.600 ;
        RECT 51.510 198.210 54.170 198.910 ;
        RECT 51.510 196.250 52.265 198.210 ;
        RECT 58.885 197.080 59.185 202.825 ;
        RECT 95.500 202.595 96.200 213.755 ;
        RECT 98.725 213.165 99.315 213.340 ;
        RECT 93.680 202.580 96.200 202.595 ;
        RECT 63.665 201.775 64.245 202.415 ;
        RECT 64.880 201.895 96.200 202.580 ;
        RECT 96.640 212.865 99.315 213.165 ;
        RECT 96.640 205.970 96.940 212.865 ;
        RECT 98.725 212.690 99.315 212.865 ;
        RECT 104.350 211.885 104.950 213.755 ;
        RECT 107.005 213.085 107.595 213.340 ;
        RECT 104.335 211.235 104.950 211.885 ;
        RECT 97.360 210.070 97.960 210.710 ;
        RECT 102.790 206.900 103.380 207.550 ;
        RECT 98.725 205.970 99.315 206.145 ;
        RECT 96.640 205.670 99.315 205.970 ;
        RECT 64.880 201.880 94.380 201.895 ;
        RECT 64.880 201.810 65.580 201.880 ;
        RECT 58.740 196.430 59.330 197.080 ;
        RECT 51.510 193.985 52.210 196.250 ;
        RECT 53.280 195.005 53.870 195.180 ;
        RECT 58.885 195.005 59.185 196.430 ;
        RECT 53.280 194.705 59.185 195.005 ;
        RECT 53.280 194.530 53.870 194.705 ;
        RECT 51.510 193.285 54.225 193.985 ;
        RECT 51.510 192.260 52.210 193.285 ;
        RECT 51.510 191.560 52.225 192.260 ;
        RECT 58.885 192.035 59.185 194.705 ;
        RECT 58.740 191.385 59.330 192.035 ;
        RECT 53.280 190.185 53.870 190.360 ;
        RECT 58.885 190.185 59.185 191.385 ;
        RECT 53.280 189.885 59.185 190.185 ;
        RECT 53.280 189.710 53.870 189.885 ;
        RECT 53.425 187.430 53.725 189.710 ;
        RECT 53.215 186.790 53.795 187.430 ;
        RECT 37.425 185.900 47.045 185.950 ;
        RECT 37.425 185.250 55.625 185.900 ;
        RECT 37.425 181.220 43.100 185.250 ;
        RECT 44.330 183.990 45.030 185.250 ;
        RECT 46.345 185.200 55.625 185.250 ;
        RECT 53.600 183.115 54.190 183.765 ;
        RECT 52.590 181.765 53.180 181.940 ;
        RECT 53.745 181.765 54.045 183.115 ;
        RECT 54.205 181.765 54.785 181.930 ;
        RECT 52.590 181.465 54.785 181.765 ;
        RECT 52.590 181.290 53.180 181.465 ;
        RECT 37.425 180.520 46.990 181.220 ;
        RECT 37.425 176.645 43.100 180.520 ;
        RECT 44.320 179.535 45.020 180.520 ;
        RECT 53.745 179.310 54.045 181.465 ;
        RECT 54.205 181.290 54.785 181.465 ;
        RECT 53.600 178.660 54.190 179.310 ;
        RECT 52.590 177.250 53.180 177.425 ;
        RECT 53.745 177.250 54.045 178.660 ;
        RECT 52.590 176.950 54.045 177.250 ;
        RECT 52.590 176.775 53.180 176.950 ;
        RECT 37.425 176.630 46.880 176.645 ;
        RECT 37.425 175.980 46.990 176.630 ;
        RECT 37.425 175.945 46.880 175.980 ;
        RECT 37.425 171.105 43.100 175.945 ;
        RECT 44.320 174.935 45.020 175.945 ;
        RECT 53.745 174.615 54.045 176.950 ;
        RECT 54.925 175.535 55.625 185.200 ;
        RECT 56.390 184.105 56.970 184.280 ;
        RECT 63.805 184.105 64.105 201.775 ;
        RECT 83.060 200.280 83.760 201.880 ;
        RECT 81.290 199.580 83.760 200.280 ;
        RECT 75.980 197.485 76.560 198.125 ;
        RECT 76.140 197.095 76.440 197.485 ;
        RECT 76.005 196.445 76.595 197.095 ;
        RECT 76.140 194.025 76.440 196.445 ;
        RECT 77.450 194.025 78.040 194.200 ;
        RECT 76.140 193.725 78.040 194.025 ;
        RECT 76.140 189.820 76.440 193.725 ;
        RECT 77.450 193.550 78.040 193.725 ;
        RECT 83.060 193.175 83.760 199.580 ;
        RECT 81.290 192.475 83.760 193.175 ;
        RECT 83.060 191.375 83.760 192.475 ;
        RECT 96.640 198.995 96.940 205.670 ;
        RECT 98.725 205.495 99.315 205.670 ;
        RECT 97.360 202.895 97.960 203.535 ;
        RECT 102.875 199.835 103.465 200.485 ;
        RECT 98.725 198.995 99.315 199.170 ;
        RECT 96.640 198.695 99.315 198.995 ;
        RECT 96.640 191.985 96.940 198.695 ;
        RECT 98.725 198.520 99.315 198.695 ;
        RECT 97.360 195.945 97.960 196.585 ;
        RECT 102.875 192.955 103.465 193.605 ;
        RECT 98.725 191.985 99.315 192.195 ;
        RECT 96.640 191.685 99.315 191.985 ;
        RECT 75.985 189.170 76.575 189.820 ;
        RECT 76.130 187.195 76.430 189.170 ;
        RECT 95.590 188.870 96.190 189.510 ;
        RECT 77.450 187.195 78.040 187.335 ;
        RECT 76.130 186.895 78.040 187.195 ;
        RECT 76.130 186.080 76.430 186.895 ;
        RECT 77.450 186.685 78.040 186.895 ;
        RECT 95.740 186.080 96.040 188.870 ;
        RECT 76.130 185.780 96.040 186.080 ;
        RECT 76.130 185.775 76.430 185.780 ;
        RECT 96.640 185.100 96.940 191.685 ;
        RECT 98.725 191.545 99.315 191.685 ;
        RECT 104.350 189.705 104.950 211.235 ;
        RECT 105.220 212.945 107.595 213.085 ;
        RECT 105.220 205.890 105.360 212.945 ;
        RECT 107.005 212.690 107.595 212.945 ;
        RECT 113.730 211.760 114.430 213.755 ;
        RECT 112.435 211.060 114.430 211.760 ;
        RECT 105.555 210.210 106.155 210.850 ;
        RECT 106.710 206.900 107.300 207.550 ;
        RECT 107.005 205.890 107.595 206.145 ;
        RECT 105.220 205.750 107.595 205.890 ;
        RECT 105.220 198.985 105.360 205.750 ;
        RECT 107.005 205.495 107.595 205.750 ;
        RECT 113.730 204.995 114.430 211.060 ;
        RECT 112.435 204.295 114.430 204.995 ;
        RECT 105.555 203.130 106.155 203.770 ;
        RECT 106.795 199.835 107.385 200.485 ;
        RECT 107.005 198.985 107.595 199.240 ;
        RECT 105.220 198.845 107.595 198.985 ;
        RECT 105.220 192.005 105.360 198.845 ;
        RECT 107.005 198.590 107.595 198.845 ;
        RECT 112.380 197.800 113.080 197.860 ;
        RECT 113.730 197.800 114.430 204.295 ;
        RECT 112.380 197.100 114.430 197.800 ;
        RECT 105.555 196.260 106.155 196.900 ;
        RECT 106.795 192.955 107.385 193.605 ;
        RECT 107.005 192.005 107.595 192.260 ;
        RECT 105.220 191.865 107.595 192.005 ;
        RECT 97.360 188.920 97.960 189.560 ;
        RECT 102.875 185.795 103.465 186.445 ;
        RECT 105.220 185.100 105.360 191.865 ;
        RECT 107.005 191.610 107.595 191.865 ;
        RECT 113.730 190.380 114.430 197.100 ;
        RECT 119.920 190.380 124.425 214.935 ;
        RECT 112.435 189.680 124.425 190.380 ;
        RECT 105.555 188.920 106.155 189.560 ;
        RECT 106.795 185.795 107.385 186.445 ;
        RECT 96.640 184.800 119.500 185.100 ;
        RECT 56.390 183.805 64.105 184.105 ;
        RECT 56.390 183.640 56.970 183.805 ;
        RECT 58.285 181.170 58.515 183.030 ;
        RECT 118.620 182.830 118.850 183.030 ;
        RECT 119.200 182.830 119.500 184.800 ;
        RECT 118.620 182.690 119.500 182.830 ;
        RECT 118.620 182.380 118.850 182.690 ;
        RECT 58.285 178.750 58.515 180.610 ;
        RECT 118.620 179.960 118.850 181.820 ;
        RECT 58.285 176.330 58.515 178.190 ;
        RECT 118.620 177.540 118.850 179.400 ;
        RECT 119.920 176.980 124.425 189.680 ;
        RECT 118.620 176.330 124.425 176.980 ;
        RECT 54.925 174.835 88.460 175.535 ;
        RECT 53.600 173.965 54.190 174.615 ;
        RECT 52.590 172.645 53.180 172.825 ;
        RECT 53.745 172.645 54.045 173.965 ;
        RECT 52.590 172.345 54.045 172.645 ;
        RECT 52.590 172.175 53.180 172.345 ;
        RECT 37.425 171.060 46.480 171.105 ;
        RECT 37.425 170.410 46.905 171.060 ;
        RECT 37.425 170.405 46.480 170.410 ;
        RECT 37.425 166.625 43.100 170.405 ;
        RECT 44.320 169.390 45.020 170.405 ;
        RECT 53.745 168.905 54.045 172.345 ;
        RECT 87.760 171.680 88.460 174.835 ;
        RECT 104.650 173.335 113.505 174.035 ;
        RECT 88.990 172.675 89.580 173.325 ;
        RECT 87.635 170.670 88.585 171.680 ;
        RECT 104.650 171.410 105.350 173.335 ;
        RECT 106.825 173.165 107.415 173.335 ;
        RECT 90.930 170.710 105.350 171.410 ;
        RECT 112.805 172.075 113.505 173.335 ;
        RECT 119.920 172.075 124.425 176.330 ;
        RECT 112.805 171.375 124.425 172.075 ;
        RECT 53.575 168.255 54.165 168.905 ;
        RECT 37.425 165.925 46.960 166.625 ;
        RECT 52.355 166.575 52.945 167.225 ;
        RECT 37.425 161.970 43.100 165.925 ;
        RECT 44.400 164.775 45.100 165.925 ;
        RECT 53.745 164.595 54.045 168.255 ;
        RECT 53.605 163.945 54.195 164.595 ;
        RECT 46.260 161.970 46.960 162.035 ;
        RECT 37.425 161.270 46.960 161.970 ;
        RECT 52.290 161.940 52.880 162.590 ;
        RECT 37.425 136.010 43.100 161.270 ;
        RECT 44.320 160.285 45.020 161.270 ;
        RECT 53.745 159.995 54.045 163.945 ;
        RECT 87.760 161.720 88.460 170.670 ;
        RECT 89.015 168.705 89.605 169.355 ;
        RECT 89.005 162.615 89.595 163.265 ;
        RECT 87.725 160.710 88.675 161.720 ;
        RECT 92.040 161.490 92.740 170.710 ;
        RECT 105.525 169.855 106.125 170.495 ;
        RECT 107.045 167.900 107.635 167.990 ;
        RECT 104.925 167.600 107.635 167.900 ;
        RECT 93.730 163.080 94.320 163.295 ;
        RECT 104.925 163.080 105.225 167.600 ;
        RECT 107.045 167.340 107.635 167.600 ;
        RECT 106.770 166.590 107.470 166.645 ;
        RECT 106.770 165.890 113.495 166.590 ;
        RECT 112.795 165.520 113.495 165.890 ;
        RECT 119.920 165.520 124.425 171.375 ;
        RECT 112.795 164.845 124.425 165.520 ;
        RECT 112.850 164.820 124.425 164.845 ;
        RECT 93.730 162.780 105.225 163.080 ;
        RECT 105.525 163.065 106.125 163.705 ;
        RECT 93.730 162.645 94.320 162.780 ;
        RECT 90.940 160.790 92.740 161.490 ;
        RECT 104.925 160.685 105.225 162.780 ;
        RECT 107.045 160.685 107.635 160.860 ;
        RECT 104.925 160.385 107.635 160.685 ;
        RECT 107.045 160.210 107.635 160.385 ;
        RECT 53.585 159.345 54.175 159.995 ;
        RECT 85.875 159.205 86.490 159.210 ;
        RECT 85.840 157.840 86.490 159.205 ;
        RECT 89.015 158.715 89.605 159.365 ;
        RECT 52.295 157.190 52.885 157.840 ;
        RECT 55.235 157.140 113.380 157.840 ;
        RECT 85.840 157.130 86.490 157.140 ;
        RECT 112.680 155.370 113.380 157.140 ;
        RECT 45.645 153.510 45.875 155.370 ;
        RECT 110.650 154.720 113.380 155.370 ;
        RECT 45.645 151.090 45.875 152.950 ;
        RECT 110.650 152.300 110.880 154.160 ;
        RECT 45.645 148.670 45.875 150.530 ;
        RECT 110.650 149.880 110.880 151.740 ;
        RECT 45.645 146.250 45.875 148.110 ;
        RECT 110.650 147.460 110.880 149.320 ;
        RECT 45.645 143.830 45.875 145.690 ;
        RECT 110.650 145.040 110.880 146.900 ;
        RECT 45.645 141.410 45.875 143.270 ;
        RECT 110.650 142.620 110.880 144.480 ;
        RECT 112.680 142.945 113.380 154.720 ;
        RECT 45.645 138.990 45.875 140.850 ;
        RECT 110.650 140.200 110.880 142.060 ;
        RECT 45.645 136.570 45.875 138.430 ;
        RECT 110.650 137.780 110.880 139.640 ;
        RECT 110.650 136.570 111.950 137.220 ;
        RECT 111.300 136.010 111.950 136.570 ;
        RECT 37.425 135.360 111.950 136.010 ;
        RECT 37.425 135.045 43.100 135.360 ;
        RECT 112.425 135.045 117.425 142.945 ;
        RECT 119.920 135.045 124.425 164.820 ;
        RECT 114.565 122.705 115.565 135.045 ;
        RECT 30.595 110.745 36.705 111.555 ;
        RECT 10.685 109.745 36.705 110.745 ;
        RECT 125.970 110.345 130.850 111.555 ;
        RECT 30.595 89.340 36.705 109.745 ;
        RECT 45.860 109.305 46.760 109.465 ;
        RECT 54.845 109.315 55.745 109.475 ;
        RECT 65.080 109.315 65.980 109.475 ;
        RECT 45.840 108.665 46.780 109.305 ;
        RECT 54.825 108.675 55.765 109.315 ;
        RECT 65.060 108.675 66.000 109.315 ;
        RECT 73.485 109.290 74.065 109.930 ;
        RECT 78.585 109.840 79.485 110.000 ;
        RECT 45.860 108.505 46.760 108.665 ;
        RECT 54.845 108.515 55.745 108.675 ;
        RECT 65.080 108.515 65.980 108.675 ;
        RECT 44.105 106.790 45.005 106.950 ;
        RECT 44.085 106.150 45.025 106.790 ;
        RECT 61.320 106.645 62.220 106.805 ;
        RECT 71.345 106.645 72.245 106.805 ;
        RECT 44.105 105.990 45.005 106.150 ;
        RECT 51.555 105.855 52.145 106.505 ;
        RECT 61.300 106.005 62.240 106.645 ;
        RECT 71.325 106.005 72.265 106.645 ;
        RECT 73.595 106.300 73.735 109.290 ;
        RECT 78.565 109.200 79.505 109.840 ;
        RECT 125.970 109.345 134.165 110.345 ;
        RECT 78.585 109.040 79.485 109.200 ;
        RECT 81.770 107.725 82.350 107.910 ;
        RECT 125.970 107.725 130.850 109.345 ;
        RECT 81.725 107.025 130.850 107.725 ;
        RECT 45.785 102.320 46.785 103.320 ;
        RECT 45.860 100.455 46.760 100.615 ;
        RECT 45.840 99.815 46.780 100.455 ;
        RECT 45.860 99.655 46.760 99.815 ;
        RECT 51.795 97.630 51.935 105.855 ;
        RECT 61.320 105.845 62.220 106.005 ;
        RECT 71.345 105.845 72.245 106.005 ;
        RECT 73.355 105.650 73.945 106.300 ;
        RECT 82.175 106.020 82.755 106.215 ;
        RECT 82.175 105.880 83.125 106.020 ;
        RECT 53.995 103.890 54.585 104.540 ;
        RECT 51.780 97.430 51.935 97.630 ;
        RECT 44.105 96.995 45.005 97.155 ;
        RECT 44.085 96.355 45.025 96.995 ;
        RECT 51.780 96.395 51.920 97.430 ;
        RECT 44.105 96.195 45.005 96.355 ;
        RECT 51.575 95.745 52.165 96.395 ;
        RECT 45.785 92.410 46.785 93.410 ;
        RECT 37.185 89.340 37.765 89.590 ;
        RECT 30.595 89.200 37.765 89.340 ;
        RECT 45.860 89.235 46.760 89.395 ;
        RECT 30.595 58.345 36.705 89.200 ;
        RECT 37.185 88.950 37.765 89.200 ;
        RECT 45.840 88.595 46.780 89.235 ;
        RECT 45.860 88.435 46.760 88.595 ;
        RECT 44.105 87.635 45.005 87.795 ;
        RECT 44.085 86.995 45.025 87.635 ;
        RECT 44.105 86.835 45.005 86.995 ;
        RECT 51.780 86.320 51.920 95.745 ;
        RECT 54.220 94.610 54.360 103.890 ;
        RECT 64.155 103.860 64.745 104.510 ;
        RECT 54.770 102.355 55.770 103.355 ;
        RECT 64.375 100.180 64.515 103.860 ;
        RECT 65.265 102.295 66.265 103.295 ;
        RECT 73.595 102.965 73.735 105.650 ;
        RECT 82.175 105.575 82.755 105.880 ;
        RECT 82.985 105.075 83.125 105.880 ;
        RECT 82.930 104.425 83.160 105.075 ;
        RECT 74.205 102.965 75.155 103.335 ;
        RECT 73.595 102.825 75.155 102.965 ;
        RECT 79.235 102.930 80.135 103.090 ;
        RECT 73.595 100.180 73.735 102.825 ;
        RECT 74.205 102.325 75.155 102.825 ;
        RECT 79.215 102.290 80.155 102.930 ;
        RECT 79.235 102.130 80.135 102.290 ;
        RECT 82.930 102.005 83.160 103.865 ;
        RECT 123.765 103.215 123.995 105.075 ;
        RECT 64.375 100.040 73.735 100.180 ;
        RECT 54.845 99.355 55.745 99.515 ;
        RECT 54.825 98.715 55.765 99.355 ;
        RECT 54.845 98.555 55.745 98.715 ;
        RECT 64.375 98.315 64.515 100.040 ;
        RECT 65.080 99.375 65.980 99.535 ;
        RECT 65.060 98.735 66.000 99.375 ;
        RECT 65.080 98.575 65.980 98.735 ;
        RECT 64.155 97.665 64.745 98.315 ;
        RECT 61.320 96.295 62.220 96.455 ;
        RECT 61.300 95.655 62.240 96.295 ;
        RECT 61.320 95.495 62.220 95.655 ;
        RECT 53.995 93.960 54.585 94.610 ;
        RECT 51.555 85.670 52.145 86.320 ;
        RECT 45.785 82.255 46.785 83.255 ;
        RECT 45.860 80.160 46.760 80.320 ;
        RECT 45.840 79.520 46.780 80.160 ;
        RECT 45.860 79.360 46.760 79.520 ;
        RECT 43.500 77.150 44.400 77.310 ;
        RECT 43.480 76.510 44.420 77.150 ;
        RECT 51.780 77.120 51.920 85.670 ;
        RECT 54.220 84.560 54.360 93.960 ;
        RECT 54.770 92.445 55.770 93.445 ;
        RECT 54.845 89.585 55.745 89.745 ;
        RECT 54.825 88.945 55.765 89.585 ;
        RECT 54.845 88.785 55.745 88.945 ;
        RECT 64.375 88.310 64.515 97.665 ;
        RECT 71.345 96.295 72.245 96.455 ;
        RECT 73.595 96.335 73.735 100.040 ;
        RECT 78.510 99.840 79.410 100.000 ;
        RECT 78.490 99.200 79.430 99.840 ;
        RECT 82.930 99.585 83.160 101.445 ;
        RECT 123.765 100.795 123.995 102.655 ;
        RECT 125.970 100.240 130.850 107.025 ;
        RECT 123.890 100.235 130.850 100.240 ;
        RECT 123.765 99.585 130.850 100.235 ;
        RECT 123.890 99.540 130.850 99.585 ;
        RECT 78.510 99.040 79.410 99.200 ;
        RECT 125.970 99.040 130.850 99.540 ;
        RECT 122.010 98.340 130.850 99.040 ;
        RECT 93.335 97.865 112.645 98.005 ;
        RECT 71.325 95.655 72.265 96.295 ;
        RECT 73.375 95.685 73.965 96.335 ;
        RECT 93.335 96.275 93.475 97.865 ;
        RECT 112.505 96.870 112.645 97.865 ;
        RECT 93.220 96.005 93.810 96.275 ;
        RECT 86.055 95.865 93.810 96.005 ;
        RECT 71.345 95.495 72.245 95.655 ;
        RECT 65.265 92.400 66.265 93.400 ;
        RECT 73.595 92.955 73.735 95.685 ;
        RECT 74.205 92.955 75.155 93.435 ;
        RECT 79.235 93.410 80.135 93.570 ;
        RECT 73.595 92.815 75.155 92.955 ;
        RECT 65.080 89.710 65.980 89.870 ;
        RECT 65.060 89.070 66.000 89.710 ;
        RECT 65.080 88.910 65.980 89.070 ;
        RECT 64.155 87.660 64.745 88.310 ;
        RECT 61.320 86.275 62.220 86.435 ;
        RECT 61.300 85.635 62.240 86.275 ;
        RECT 61.320 85.475 62.220 85.635 ;
        RECT 53.995 83.910 54.585 84.560 ;
        RECT 54.210 80.970 54.350 83.910 ;
        RECT 54.770 82.430 55.770 83.430 ;
        RECT 64.380 80.970 64.520 87.660 ;
        RECT 71.345 86.435 72.245 86.595 ;
        RECT 73.595 86.575 73.735 92.815 ;
        RECT 74.205 92.425 75.155 92.815 ;
        RECT 79.215 92.770 80.155 93.410 ;
        RECT 79.235 92.610 80.135 92.770 ;
        RECT 78.510 90.010 79.410 90.170 ;
        RECT 78.490 89.370 79.430 90.010 ;
        RECT 78.510 89.210 79.410 89.370 ;
        RECT 71.325 85.795 72.265 86.435 ;
        RECT 73.315 85.925 73.905 86.575 ;
        RECT 71.345 85.635 72.245 85.795 ;
        RECT 73.595 84.670 73.735 85.925 ;
        RECT 73.580 84.530 73.735 84.670 ;
        RECT 65.265 82.545 66.265 83.545 ;
        RECT 54.210 80.830 64.520 80.970 ;
        RECT 54.210 79.140 54.350 80.830 ;
        RECT 54.845 80.150 55.745 80.310 ;
        RECT 54.825 79.510 55.765 80.150 ;
        RECT 54.845 79.350 55.745 79.510 ;
        RECT 53.995 78.490 54.585 79.140 ;
        RECT 64.380 79.045 64.520 80.830 ;
        RECT 65.080 80.195 65.980 80.355 ;
        RECT 65.060 79.555 66.000 80.195 ;
        RECT 65.080 79.395 65.980 79.555 ;
        RECT 64.155 78.395 64.745 79.045 ;
        RECT 61.320 77.340 62.220 77.500 ;
        RECT 51.575 76.855 52.165 77.120 ;
        RECT 52.350 76.855 52.930 77.105 ;
        RECT 51.575 76.715 52.930 76.855 ;
        RECT 43.500 76.350 44.400 76.510 ;
        RECT 51.575 76.470 52.165 76.715 ;
        RECT 52.350 76.465 52.930 76.715 ;
        RECT 61.300 76.700 62.240 77.340 ;
        RECT 71.345 77.110 72.245 77.270 ;
        RECT 61.320 76.540 62.220 76.700 ;
        RECT 71.325 76.470 72.265 77.110 ;
        RECT 73.595 76.875 73.735 84.530 ;
        RECT 74.310 82.695 75.310 83.695 ;
        RECT 79.200 83.055 80.100 83.215 ;
        RECT 79.180 82.415 80.120 83.055 ;
        RECT 79.200 82.255 80.100 82.415 ;
        RECT 78.670 79.885 79.570 80.045 ;
        RECT 78.650 79.245 79.590 79.885 ;
        RECT 78.670 79.085 79.570 79.245 ;
        RECT 86.055 77.260 86.195 95.865 ;
        RECT 93.220 95.625 93.810 95.865 ;
        RECT 96.455 95.620 97.455 96.620 ;
        RECT 97.960 96.245 98.860 96.405 ;
        RECT 97.940 95.605 98.880 96.245 ;
        RECT 112.255 96.220 112.845 96.870 ;
        RECT 114.785 95.620 115.785 96.620 ;
        RECT 116.290 96.245 117.190 96.405 ;
        RECT 116.270 95.605 117.210 96.245 ;
        RECT 97.960 95.445 98.860 95.605 ;
        RECT 116.290 95.445 117.190 95.605 ;
        RECT 96.030 94.995 96.930 95.155 ;
        RECT 114.360 94.995 115.260 95.155 ;
        RECT 94.550 93.895 95.550 94.895 ;
        RECT 96.010 94.355 96.950 94.995 ;
        RECT 96.030 94.195 96.930 94.355 ;
        RECT 93.520 92.330 94.520 93.330 ;
        RECT 94.980 93.325 95.880 93.485 ;
        RECT 94.960 92.685 95.900 93.325 ;
        RECT 104.585 93.210 105.585 94.210 ;
        RECT 112.880 93.895 113.880 94.895 ;
        RECT 114.340 94.355 115.280 94.995 ;
        RECT 114.360 94.195 115.260 94.355 ;
        RECT 94.980 92.525 95.880 92.685 ;
        RECT 111.850 92.330 112.850 93.330 ;
        RECT 113.310 93.325 114.210 93.485 ;
        RECT 113.290 92.685 114.230 93.325 ;
        RECT 113.310 92.525 114.210 92.685 ;
        RECT 89.665 90.930 90.565 91.090 ;
        RECT 89.645 90.290 90.585 90.930 ;
        RECT 91.170 90.825 92.170 91.825 ;
        RECT 92.865 91.745 93.765 91.905 ;
        RECT 92.845 91.105 93.785 91.745 ;
        RECT 92.865 90.945 93.765 91.105 ;
        RECT 107.995 90.930 108.895 91.090 ;
        RECT 107.975 90.290 108.915 90.930 ;
        RECT 109.500 90.825 110.500 91.825 ;
        RECT 111.195 91.745 112.095 91.905 ;
        RECT 111.175 91.105 112.115 91.745 ;
        RECT 111.195 90.945 112.095 91.105 ;
        RECT 89.665 90.130 90.565 90.290 ;
        RECT 107.995 90.130 108.895 90.290 ;
        RECT 87.955 88.665 88.955 89.665 ;
        RECT 89.665 88.570 90.565 88.730 ;
        RECT 106.285 88.685 107.285 89.685 ;
        RECT 125.970 89.640 130.850 98.340 ;
        RECT 121.875 88.940 130.850 89.640 ;
        RECT 107.995 88.570 108.895 88.730 ;
        RECT 89.645 87.930 90.585 88.570 ;
        RECT 107.975 87.930 108.915 88.570 ;
        RECT 89.665 87.770 90.565 87.930 ;
        RECT 107.995 87.770 108.895 87.930 ;
        RECT 90.490 86.285 91.490 87.285 ;
        RECT 92.000 87.105 92.900 87.265 ;
        RECT 91.980 86.465 92.920 87.105 ;
        RECT 92.000 86.305 92.900 86.465 ;
        RECT 108.820 86.285 109.820 87.285 ;
        RECT 110.330 87.105 111.230 87.265 ;
        RECT 110.310 86.465 111.250 87.105 ;
        RECT 110.330 86.305 111.230 86.465 ;
        RECT 92.565 84.860 93.565 85.860 ;
        RECT 94.105 85.585 95.005 85.745 ;
        RECT 94.085 84.945 95.025 85.585 ;
        RECT 94.105 84.785 95.005 84.945 ;
        RECT 110.895 84.860 111.895 85.860 ;
        RECT 112.435 85.585 113.335 85.745 ;
        RECT 112.415 84.945 113.355 85.585 ;
        RECT 112.435 84.785 113.335 84.945 ;
        RECT 92.565 82.915 93.565 83.915 ;
        RECT 94.310 83.760 95.210 83.920 ;
        RECT 94.290 83.120 95.230 83.760 ;
        RECT 94.310 82.960 95.210 83.120 ;
        RECT 110.895 82.915 111.895 83.915 ;
        RECT 112.640 83.760 113.540 83.920 ;
        RECT 112.620 83.120 113.560 83.760 ;
        RECT 112.640 82.960 113.540 83.120 ;
        RECT 94.835 81.375 95.835 82.375 ;
        RECT 96.390 82.300 97.290 82.460 ;
        RECT 96.370 81.660 97.310 82.300 ;
        RECT 96.390 81.500 97.290 81.660 ;
        RECT 97.990 81.375 98.990 82.375 ;
        RECT 113.165 81.375 114.165 82.375 ;
        RECT 114.720 82.300 115.620 82.460 ;
        RECT 114.700 81.660 115.640 82.300 ;
        RECT 114.720 81.500 115.620 81.660 ;
        RECT 116.320 81.375 117.320 82.375 ;
        RECT 93.085 79.025 111.925 79.165 ;
        RECT 93.085 77.890 93.225 79.025 ;
        RECT 92.910 77.260 93.500 77.890 ;
        RECT 96.215 77.330 97.215 78.330 ;
        RECT 97.670 77.955 98.570 78.115 ;
        RECT 97.650 77.315 98.590 77.955 ;
        RECT 111.785 77.515 111.925 79.025 ;
        RECT 86.055 77.240 93.500 77.260 ;
        RECT 86.055 77.120 93.225 77.240 ;
        RECT 97.670 77.155 98.570 77.315 ;
        RECT 71.345 76.310 72.245 76.470 ;
        RECT 73.335 76.225 73.925 76.875 ;
        RECT 45.785 73.250 46.785 74.250 ;
        RECT 54.770 73.225 55.770 74.225 ;
        RECT 65.265 73.370 66.265 74.370 ;
        RECT 73.905 73.070 74.905 74.070 ;
        RECT 79.330 73.535 80.230 73.695 ;
        RECT 79.310 72.895 80.250 73.535 ;
        RECT 79.330 72.735 80.230 72.895 ;
        RECT 51.545 72.155 52.445 72.315 ;
        RECT 51.525 71.515 52.465 72.155 ;
        RECT 51.545 71.355 52.445 71.515 ;
        RECT 58.270 69.570 58.850 70.210 ;
        RECT 58.455 68.865 58.595 69.570 ;
        RECT 74.360 69.400 74.940 69.650 ;
        RECT 75.620 69.400 76.210 69.655 ;
        RECT 63.540 69.185 64.440 69.345 ;
        RECT 74.360 69.260 76.210 69.400 ;
        RECT 58.230 68.215 58.820 68.865 ;
        RECT 63.520 68.545 64.460 69.185 ;
        RECT 74.360 69.010 74.940 69.260 ;
        RECT 75.620 69.005 76.210 69.260 ;
        RECT 63.540 68.385 64.440 68.545 ;
        RECT 51.380 66.050 52.380 67.050 ;
        RECT 51.545 65.615 52.445 65.775 ;
        RECT 51.525 64.975 52.465 65.615 ;
        RECT 51.545 64.815 52.445 64.975 ;
        RECT 58.470 63.530 58.610 68.215 ;
        RECT 63.540 67.365 64.440 67.525 ;
        RECT 63.520 66.725 64.460 67.365 ;
        RECT 75.845 67.140 75.985 69.005 ;
        RECT 63.540 66.565 64.440 66.725 ;
        RECT 75.620 66.490 76.210 67.140 ;
        RECT 63.540 65.545 64.440 65.705 ;
        RECT 63.520 64.905 64.460 65.545 ;
        RECT 63.540 64.745 64.440 64.905 ;
        RECT 75.845 64.535 75.985 66.490 ;
        RECT 63.550 63.730 64.450 63.890 ;
        RECT 75.620 63.885 76.210 64.535 ;
        RECT 58.250 62.880 58.840 63.530 ;
        RECT 63.530 63.090 64.470 63.730 ;
        RECT 63.550 62.930 64.450 63.090 ;
        RECT 47.830 59.945 48.410 60.175 ;
        RECT 45.140 59.805 48.410 59.945 ;
        RECT 30.595 58.330 37.700 58.345 ;
        RECT 30.595 57.690 37.990 58.330 ;
        RECT 30.595 57.645 37.700 57.690 ;
        RECT 30.595 47.670 36.705 57.645 ;
        RECT 30.595 46.970 37.990 47.670 ;
        RECT 30.595 46.115 36.705 46.970 ;
        RECT 37.220 46.115 38.530 46.460 ;
        RECT 30.595 45.415 38.530 46.115 ;
        RECT 43.635 45.690 44.535 45.850 ;
        RECT 30.595 39.535 36.705 45.415 ;
        RECT 37.220 45.090 38.530 45.415 ;
        RECT 43.615 45.050 44.555 45.690 ;
        RECT 43.635 44.890 44.535 45.050 ;
        RECT 45.140 43.315 45.280 59.805 ;
        RECT 47.830 59.535 48.410 59.805 ;
        RECT 51.380 59.360 52.380 60.360 ;
        RECT 51.545 58.920 52.445 59.080 ;
        RECT 51.525 58.280 52.465 58.920 ;
        RECT 51.545 58.120 52.445 58.280 ;
        RECT 58.455 55.045 58.595 62.880 ;
        RECT 63.550 61.905 64.450 62.065 ;
        RECT 75.845 62.005 75.985 63.885 ;
        RECT 63.530 61.265 64.470 61.905 ;
        RECT 75.620 61.355 76.210 62.005 ;
        RECT 63.550 61.105 64.450 61.265 ;
        RECT 63.550 60.080 64.450 60.240 ;
        RECT 63.530 59.440 64.470 60.080 ;
        RECT 63.550 59.280 64.450 59.440 ;
        RECT 75.845 59.360 75.985 61.355 ;
        RECT 75.620 58.710 76.210 59.360 ;
        RECT 63.540 58.270 64.440 58.430 ;
        RECT 63.520 57.630 64.460 58.270 ;
        RECT 63.540 57.470 64.440 57.630 ;
        RECT 75.845 56.885 75.985 58.710 ;
        RECT 61.245 56.445 62.145 56.605 ;
        RECT 63.550 56.445 64.450 56.605 ;
        RECT 61.225 55.805 62.165 56.445 ;
        RECT 63.530 55.805 64.470 56.445 ;
        RECT 75.620 56.235 76.210 56.885 ;
        RECT 73.040 55.960 73.620 56.225 ;
        RECT 74.295 55.960 74.885 56.215 ;
        RECT 73.040 55.820 74.885 55.960 ;
        RECT 61.245 55.645 62.145 55.805 ;
        RECT 63.550 55.645 64.450 55.805 ;
        RECT 73.040 55.585 73.620 55.820 ;
        RECT 74.295 55.565 74.885 55.820 ;
        RECT 86.055 55.490 86.195 77.120 ;
        RECT 111.560 76.865 112.150 77.515 ;
        RECT 114.815 77.085 115.815 78.085 ;
        RECT 116.320 77.710 117.220 77.870 ;
        RECT 116.300 77.070 117.240 77.710 ;
        RECT 116.320 76.910 117.220 77.070 ;
        RECT 95.740 76.705 96.640 76.865 ;
        RECT 94.260 75.605 95.260 76.605 ;
        RECT 95.720 76.065 96.660 76.705 ;
        RECT 114.390 76.460 115.290 76.620 ;
        RECT 95.740 75.905 96.640 76.065 ;
        RECT 112.910 75.360 113.910 76.360 ;
        RECT 114.370 75.820 115.310 76.460 ;
        RECT 114.390 75.660 115.290 75.820 ;
        RECT 93.230 74.040 94.230 75.040 ;
        RECT 94.690 75.035 95.590 75.195 ;
        RECT 94.670 74.395 95.610 75.035 ;
        RECT 94.690 74.235 95.590 74.395 ;
        RECT 111.880 73.795 112.880 74.795 ;
        RECT 113.340 74.790 114.240 74.950 ;
        RECT 113.320 74.150 114.260 74.790 ;
        RECT 113.340 73.990 114.240 74.150 ;
        RECT 89.375 72.640 90.275 72.800 ;
        RECT 89.355 72.000 90.295 72.640 ;
        RECT 90.880 72.535 91.880 73.535 ;
        RECT 92.575 73.455 93.475 73.615 ;
        RECT 92.555 72.815 93.495 73.455 ;
        RECT 92.575 72.655 93.475 72.815 ;
        RECT 108.025 72.395 108.925 72.555 ;
        RECT 89.375 71.840 90.275 72.000 ;
        RECT 108.005 71.755 108.945 72.395 ;
        RECT 109.530 72.290 110.530 73.290 ;
        RECT 111.225 73.210 112.125 73.370 ;
        RECT 111.205 72.570 112.145 73.210 ;
        RECT 111.225 72.410 112.125 72.570 ;
        RECT 108.025 71.595 108.925 71.755 ;
        RECT 87.665 70.395 88.665 71.395 ;
        RECT 89.375 70.280 90.275 70.440 ;
        RECT 89.355 69.640 90.295 70.280 ;
        RECT 106.315 70.165 107.315 71.165 ;
        RECT 125.970 71.035 130.850 88.940 ;
        RECT 122.160 70.335 130.850 71.035 ;
        RECT 108.025 70.035 108.925 70.195 ;
        RECT 89.375 69.480 90.275 69.640 ;
        RECT 108.005 69.395 108.945 70.035 ;
        RECT 108.025 69.235 108.925 69.395 ;
        RECT 90.200 67.995 91.200 68.995 ;
        RECT 91.710 68.815 92.610 68.975 ;
        RECT 91.690 68.175 92.630 68.815 ;
        RECT 91.710 68.015 92.610 68.175 ;
        RECT 108.850 67.750 109.850 68.750 ;
        RECT 110.360 68.570 111.260 68.730 ;
        RECT 110.340 67.930 111.280 68.570 ;
        RECT 110.360 67.770 111.260 67.930 ;
        RECT 92.275 66.570 93.275 67.570 ;
        RECT 93.815 67.295 94.715 67.455 ;
        RECT 93.795 66.655 94.735 67.295 ;
        RECT 93.815 66.495 94.715 66.655 ;
        RECT 110.925 66.325 111.925 67.325 ;
        RECT 112.465 67.050 113.365 67.210 ;
        RECT 112.445 66.410 113.385 67.050 ;
        RECT 112.465 66.250 113.365 66.410 ;
        RECT 92.275 64.625 93.275 65.625 ;
        RECT 94.020 65.470 94.920 65.630 ;
        RECT 94.000 64.830 94.940 65.470 ;
        RECT 104.060 65.280 104.650 65.655 ;
        RECT 94.020 64.670 94.920 64.830 ;
        RECT 94.545 63.085 95.545 64.085 ;
        RECT 96.100 64.010 97.000 64.170 ;
        RECT 96.080 63.370 97.020 64.010 ;
        RECT 96.100 63.210 97.000 63.370 ;
        RECT 97.700 63.085 98.700 64.085 ;
        RECT 104.005 61.190 104.705 65.280 ;
        RECT 110.925 64.380 111.925 65.380 ;
        RECT 112.670 65.225 113.570 65.385 ;
        RECT 112.650 64.585 113.590 65.225 ;
        RECT 112.670 64.425 113.570 64.585 ;
        RECT 113.195 62.840 114.195 63.840 ;
        RECT 114.750 63.765 115.650 63.925 ;
        RECT 114.730 63.125 115.670 63.765 ;
        RECT 114.750 62.965 115.650 63.125 ;
        RECT 116.350 62.840 117.350 63.840 ;
        RECT 125.970 61.190 130.850 70.335 ;
        RECT 104.005 60.490 130.850 61.190 ;
        RECT 104.035 59.820 104.735 60.490 ;
        RECT 75.755 55.350 86.195 55.490 ;
        RECT 101.550 59.120 104.735 59.820 ;
        RECT 58.230 54.395 58.820 55.045 ;
        RECT 75.755 55.010 75.895 55.350 ;
        RECT 60.330 54.870 75.895 55.010 ;
        RECT 51.380 52.695 52.380 53.695 ;
        RECT 51.470 51.990 52.370 52.150 ;
        RECT 51.450 51.350 52.390 51.990 ;
        RECT 51.470 51.190 52.370 51.350 ;
        RECT 58.470 49.475 58.610 54.395 ;
        RECT 60.330 52.860 60.470 54.870 ;
        RECT 101.550 54.225 102.250 59.120 ;
        RECT 107.015 58.135 107.915 58.295 ;
        RECT 106.995 57.495 107.935 58.135 ;
        RECT 107.015 57.335 107.915 57.495 ;
        RECT 108.550 57.205 109.550 58.205 ;
        RECT 110.020 58.135 110.920 58.295 ;
        RECT 110.000 57.495 110.940 58.135 ;
        RECT 110.020 57.335 110.920 57.495 ;
        RECT 111.550 57.205 112.550 58.205 ;
        RECT 113.990 58.135 114.890 58.295 ;
        RECT 113.970 57.495 114.910 58.135 ;
        RECT 113.990 57.335 114.890 57.495 ;
        RECT 106.300 55.795 107.300 56.795 ;
        RECT 71.800 53.525 102.250 54.225 ;
        RECT 105.965 54.120 106.965 55.120 ;
        RECT 107.570 55.060 108.470 55.220 ;
        RECT 107.550 54.420 108.490 55.060 ;
        RECT 107.570 54.260 108.470 54.420 ;
        RECT 59.980 51.850 60.930 52.860 ;
        RECT 63.775 52.480 64.675 52.640 ;
        RECT 60.385 50.300 60.525 51.850 ;
        RECT 63.755 51.840 64.695 52.480 ;
        RECT 73.040 52.180 73.620 52.475 ;
        RECT 74.660 52.180 75.250 52.435 ;
        RECT 73.040 52.040 75.250 52.180 ;
        RECT 61.395 50.805 62.395 51.805 ;
        RECT 63.775 51.680 64.675 51.840 ;
        RECT 73.040 51.835 73.620 52.040 ;
        RECT 74.660 51.785 75.250 52.040 ;
        RECT 75.565 52.035 76.265 53.525 ;
        RECT 106.530 52.885 107.430 53.045 ;
        RECT 106.510 52.245 107.450 52.885 ;
        RECT 106.530 52.085 107.430 52.245 ;
        RECT 75.505 51.755 76.265 52.035 ;
        RECT 75.505 51.615 76.380 51.755 ;
        RECT 125.970 51.745 130.850 60.490 ;
        RECT 75.505 51.335 76.265 51.615 ;
        RECT 63.775 50.660 64.675 50.820 ;
        RECT 60.090 49.660 60.670 50.300 ;
        RECT 63.755 50.020 64.695 50.660 ;
        RECT 58.250 48.825 58.840 49.475 ;
        RECT 61.395 48.920 62.395 49.920 ;
        RECT 63.775 49.860 64.675 50.020 ;
        RECT 72.930 49.920 73.930 50.920 ;
        RECT 75.770 49.445 75.910 51.335 ;
        RECT 105.965 50.500 106.965 51.500 ;
        RECT 121.800 51.045 130.850 51.745 ;
        RECT 106.530 49.605 107.430 49.765 ;
        RECT 63.775 48.840 64.675 49.000 ;
        RECT 63.755 48.200 64.695 48.840 ;
        RECT 75.545 48.795 76.135 49.445 ;
        RECT 106.510 48.965 107.450 49.605 ;
        RECT 106.530 48.805 107.430 48.965 ;
        RECT 61.395 47.095 62.395 48.095 ;
        RECT 63.775 48.040 64.675 48.200 ;
        RECT 72.870 47.350 73.870 48.350 ;
        RECT 51.380 46.070 52.380 47.070 ;
        RECT 63.785 47.020 64.685 47.180 ;
        RECT 63.765 46.380 64.705 47.020 ;
        RECT 75.765 46.890 75.905 48.795 ;
        RECT 63.785 46.220 64.685 46.380 ;
        RECT 75.540 46.240 76.130 46.890 ;
        RECT 105.965 46.750 106.965 47.750 ;
        RECT 107.570 47.565 108.470 47.725 ;
        RECT 107.550 46.925 108.490 47.565 ;
        RECT 107.570 46.765 108.470 46.925 ;
        RECT 48.210 45.685 49.110 45.845 ;
        RECT 48.190 45.045 49.130 45.685 ;
        RECT 61.395 45.220 62.395 46.220 ;
        RECT 63.785 45.200 64.685 45.360 ;
        RECT 48.210 44.885 49.110 45.045 ;
        RECT 63.765 44.560 64.705 45.200 ;
        RECT 72.980 44.845 73.980 45.845 ;
        RECT 63.785 44.400 64.685 44.560 ;
        RECT 46.710 43.545 47.610 43.705 ;
        RECT 44.950 42.665 45.540 43.315 ;
        RECT 46.690 42.905 47.630 43.545 ;
        RECT 61.395 43.400 62.395 44.400 ;
        RECT 75.805 44.325 75.945 46.240 ;
        RECT 106.640 45.145 107.640 46.145 ;
        RECT 107.570 44.435 108.470 44.595 ;
        RECT 75.580 43.675 76.170 44.325 ;
        RECT 107.550 43.795 108.490 44.435 ;
        RECT 63.785 43.375 64.685 43.535 ;
        RECT 46.710 42.745 47.610 42.905 ;
        RECT 39.305 39.840 40.305 40.840 ;
        RECT 37.220 39.535 38.530 39.730 ;
        RECT 30.595 38.835 38.530 39.535 ;
        RECT 43.655 39.030 44.555 39.190 ;
        RECT 30.595 33.040 36.705 38.835 ;
        RECT 37.220 38.360 38.530 38.835 ;
        RECT 43.635 38.390 44.575 39.030 ;
        RECT 43.655 38.230 44.555 38.390 ;
        RECT 45.140 37.240 45.280 42.665 ;
        RECT 55.010 42.250 55.600 42.900 ;
        RECT 63.765 42.735 64.705 43.375 ;
        RECT 48.115 39.850 49.115 40.850 ;
        RECT 48.210 39.055 49.110 39.215 ;
        RECT 48.190 38.415 49.130 39.055 ;
        RECT 48.210 38.255 49.110 38.415 ;
        RECT 55.250 37.240 55.390 42.250 ;
        RECT 61.395 41.660 62.395 42.660 ;
        RECT 63.785 42.575 64.685 42.735 ;
        RECT 72.980 42.235 73.980 43.235 ;
        RECT 75.780 41.765 75.920 43.675 ;
        RECT 107.570 43.635 108.470 43.795 ;
        RECT 109.050 43.655 110.050 44.655 ;
        RECT 110.470 44.410 111.370 44.570 ;
        RECT 110.450 43.770 111.390 44.410 ;
        RECT 110.470 43.610 111.370 43.770 ;
        RECT 111.780 43.695 112.780 44.695 ;
        RECT 113.990 44.665 114.890 44.825 ;
        RECT 113.970 44.025 114.910 44.665 ;
        RECT 125.970 44.645 130.850 51.045 ;
        RECT 125.695 44.595 130.850 44.645 ;
        RECT 113.990 43.865 114.890 44.025 ;
        RECT 125.330 43.955 130.850 44.595 ;
        RECT 125.695 43.945 130.850 43.955 ;
        RECT 63.775 41.565 64.675 41.725 ;
        RECT 63.755 40.925 64.695 41.565 ;
        RECT 75.555 41.115 76.145 41.765 ;
        RECT 97.175 41.135 98.175 42.135 ;
        RECT 112.735 41.605 113.325 42.255 ;
        RECT 61.395 39.825 62.395 40.825 ;
        RECT 63.775 40.765 64.675 40.925 ;
        RECT 63.785 39.740 64.685 39.900 ;
        RECT 72.980 39.750 73.980 40.750 ;
        RECT 63.765 39.100 64.705 39.740 ;
        RECT 63.785 38.940 64.685 39.100 ;
        RECT 73.075 38.715 73.655 38.885 ;
        RECT 70.045 38.415 74.670 38.715 ;
        RECT 45.140 37.095 45.285 37.240 ;
        RECT 55.250 37.095 55.395 37.240 ;
        RECT 45.145 36.610 45.285 37.095 ;
        RECT 44.920 35.960 45.510 36.610 ;
        RECT 46.710 36.580 47.610 36.740 ;
        RECT 37.220 33.040 38.530 33.635 ;
        RECT 38.955 33.135 39.955 34.135 ;
        RECT 30.595 32.340 38.530 33.040 ;
        RECT 43.615 32.915 44.515 33.075 ;
        RECT 30.595 26.815 36.705 32.340 ;
        RECT 37.220 32.265 38.530 32.340 ;
        RECT 43.595 32.275 44.535 32.915 ;
        RECT 43.615 32.115 44.515 32.275 ;
        RECT 45.145 30.520 45.285 35.960 ;
        RECT 46.690 35.940 47.630 36.580 ;
        RECT 55.255 36.565 55.395 37.095 ;
        RECT 57.670 36.990 58.570 37.150 ;
        RECT 46.710 35.780 47.610 35.940 ;
        RECT 55.030 35.915 55.620 36.565 ;
        RECT 57.650 36.350 58.590 36.990 ;
        RECT 57.670 36.190 58.570 36.350 ;
        RECT 48.100 33.145 49.100 34.145 ;
        RECT 49.400 32.895 50.300 33.055 ;
        RECT 49.380 32.255 50.320 32.895 ;
        RECT 49.400 32.095 50.300 32.255 ;
        RECT 55.255 30.540 55.395 35.915 ;
        RECT 58.955 35.615 59.955 36.615 ;
        RECT 66.570 34.855 67.160 34.915 ;
        RECT 66.570 34.265 67.300 34.855 ;
        RECT 58.955 32.570 59.955 33.570 ;
        RECT 44.920 29.870 45.510 30.520 ;
        RECT 46.710 30.295 47.610 30.455 ;
        RECT 37.390 26.815 38.700 27.265 ;
        RECT 38.955 27.020 39.955 28.020 ;
        RECT 30.595 26.115 38.700 26.815 ;
        RECT 43.655 26.490 44.555 26.650 ;
        RECT 30.595 18.230 36.705 26.115 ;
        RECT 37.390 25.895 38.700 26.115 ;
        RECT 43.635 25.850 44.575 26.490 ;
        RECT 43.655 25.690 44.555 25.850 ;
        RECT 45.145 24.045 45.285 29.870 ;
        RECT 46.690 29.655 47.630 30.295 ;
        RECT 55.030 29.890 55.620 30.540 ;
        RECT 46.710 29.495 47.610 29.655 ;
        RECT 48.135 27.050 49.135 28.050 ;
        RECT 49.400 26.490 50.300 26.650 ;
        RECT 49.380 25.850 50.320 26.490 ;
        RECT 49.400 25.690 50.300 25.850 ;
        RECT 46.710 24.220 47.610 24.380 ;
        RECT 44.920 23.395 45.510 24.045 ;
        RECT 46.690 23.580 47.630 24.220 ;
        RECT 55.255 24.195 55.395 29.890 ;
        RECT 56.880 27.580 63.715 28.230 ;
        RECT 46.710 23.420 47.610 23.580 ;
        RECT 55.030 23.545 55.620 24.195 ;
        RECT 37.965 20.625 38.965 21.625 ;
        RECT 45.145 19.160 45.285 23.395 ;
        RECT 48.090 20.645 49.090 21.645 ;
        RECT 55.255 19.160 55.395 23.545 ;
        RECT 45.145 19.020 55.395 19.160 ;
        RECT 56.880 18.230 57.530 27.580 ;
        RECT 63.485 25.160 63.715 27.020 ;
        RECT 63.485 22.740 63.715 24.600 ;
        RECT 30.595 17.580 57.530 18.230 ;
        RECT 30.595 11.765 36.705 17.580 ;
        RECT 66.600 17.030 67.300 34.265 ;
        RECT 70.045 33.365 70.345 38.415 ;
        RECT 73.075 38.245 73.655 38.415 ;
        RECT 74.370 37.505 74.670 38.415 ;
        RECT 75.725 38.085 75.865 41.115 ;
        RECT 76.030 38.085 76.620 38.340 ;
        RECT 75.725 37.945 76.620 38.085 ;
        RECT 76.030 37.690 76.620 37.945 ;
        RECT 72.820 35.970 73.770 36.980 ;
        RECT 74.305 36.865 74.885 37.505 ;
        RECT 70.750 35.075 71.650 35.235 ;
        RECT 70.730 34.435 71.670 35.075 ;
        RECT 70.750 34.275 71.650 34.435 ;
        RECT 73.285 33.365 73.875 33.550 ;
        RECT 70.045 33.065 73.875 33.365 ;
        RECT 73.285 32.900 73.875 33.065 ;
        RECT 57.325 11.750 67.325 17.030 ;
        RECT 80.555 16.845 81.255 35.105 ;
        RECT 88.550 26.370 88.780 28.230 ;
        RECT 88.550 23.950 88.780 25.810 ;
        RECT 88.550 22.740 89.760 23.390 ;
        RECT 89.110 19.600 89.760 22.740 ;
        RECT 97.325 19.775 98.025 41.135 ;
        RECT 112.960 40.775 113.100 41.605 ;
        RECT 112.660 40.135 113.240 40.775 ;
        RECT 97.175 19.600 98.175 19.775 ;
        RECT 89.110 18.950 98.175 19.600 ;
        RECT 89.110 17.015 89.760 18.950 ;
        RECT 97.175 18.775 98.175 18.950 ;
        RECT 71.265 11.770 81.265 16.845 ;
        RECT 88.230 11.775 98.230 17.015 ;
        RECT 65.355 6.325 66.355 11.750 ;
        RECT 79.715 8.415 80.715 11.770 ;
        RECT 96.905 10.690 97.905 11.775 ;
        RECT 125.970 11.765 130.850 43.945 ;
        RECT 96.905 9.690 155.680 10.690 ;
        RECT 154.565 8.945 155.680 9.690 ;
        RECT 154.565 8.895 155.660 8.945 ;
        RECT 79.715 7.415 135.345 8.415 ;
        RECT 65.355 5.325 113.235 6.325 ;
      LAYER via ;
        RECT 59.855 218.620 60.755 219.520 ;
        RECT 10.715 213.705 11.615 214.605 ;
        RECT 127.580 214.985 128.480 215.885 ;
        RECT 53.270 205.795 53.850 206.375 ;
        RECT 63.845 206.725 64.425 207.305 ;
        RECT 92.930 206.725 93.510 207.305 ;
        RECT 63.665 202.920 64.245 203.500 ;
        RECT 92.930 202.940 93.510 203.520 ;
        RECT 53.230 200.985 53.810 201.565 ;
        RECT 63.665 201.805 64.245 202.385 ;
        RECT 97.370 210.100 97.950 210.680 ;
        RECT 102.795 206.935 103.375 207.515 ;
        RECT 53.215 186.820 53.795 187.400 ;
        RECT 54.205 181.320 54.785 181.900 ;
        RECT 56.390 183.670 56.970 184.250 ;
        RECT 75.980 197.515 76.560 198.095 ;
        RECT 97.370 202.925 97.950 203.505 ;
        RECT 102.880 199.870 103.460 200.450 ;
        RECT 97.370 195.975 97.950 196.555 ;
        RECT 102.880 192.990 103.460 193.570 ;
        RECT 95.600 188.900 96.180 189.480 ;
        RECT 105.565 210.240 106.145 210.820 ;
        RECT 106.715 206.935 107.295 207.515 ;
        RECT 105.565 203.160 106.145 203.740 ;
        RECT 106.800 199.870 107.380 200.450 ;
        RECT 105.565 196.290 106.145 196.870 ;
        RECT 106.800 192.990 107.380 193.570 ;
        RECT 97.370 188.950 97.950 189.530 ;
        RECT 102.880 185.830 103.460 186.410 ;
        RECT 105.565 188.950 106.145 189.530 ;
        RECT 106.800 185.830 107.380 186.410 ;
        RECT 88.995 172.710 89.575 173.290 ;
        RECT 52.360 166.610 52.940 167.190 ;
        RECT 52.295 161.975 52.875 162.555 ;
        RECT 89.020 168.740 89.600 169.320 ;
        RECT 89.010 162.650 89.590 163.230 ;
        RECT 105.535 169.885 106.115 170.465 ;
        RECT 93.735 162.680 94.315 163.260 ;
        RECT 105.535 163.095 106.115 163.675 ;
        RECT 85.875 158.595 86.455 159.175 ;
        RECT 89.020 158.750 89.600 159.330 ;
        RECT 52.300 157.225 52.880 157.805 ;
        RECT 55.235 157.200 55.815 157.780 ;
        RECT 114.615 122.705 115.515 123.605 ;
        RECT 10.715 109.795 11.615 110.695 ;
        RECT 45.860 108.535 46.760 109.435 ;
        RECT 54.845 108.545 55.745 109.445 ;
        RECT 65.080 108.545 65.980 109.445 ;
        RECT 73.485 109.320 74.065 109.900 ;
        RECT 44.105 106.020 45.005 106.920 ;
        RECT 61.320 105.875 62.220 106.775 ;
        RECT 45.835 102.370 46.735 103.270 ;
        RECT 45.860 99.685 46.760 100.585 ;
        RECT 71.345 105.875 72.245 106.775 ;
        RECT 78.585 109.070 79.485 109.970 ;
        RECT 133.235 109.395 134.135 110.295 ;
        RECT 81.770 107.300 82.350 107.880 ;
        RECT 44.105 96.225 45.005 97.125 ;
        RECT 45.835 92.460 46.735 93.360 ;
        RECT 37.185 88.980 37.765 89.560 ;
        RECT 45.860 88.465 46.760 89.365 ;
        RECT 44.105 86.865 45.005 87.765 ;
        RECT 54.820 102.405 55.720 103.305 ;
        RECT 65.315 102.345 66.215 103.245 ;
        RECT 82.175 105.605 82.755 106.185 ;
        RECT 79.235 102.160 80.135 103.060 ;
        RECT 54.845 98.585 55.745 99.485 ;
        RECT 65.080 98.605 65.980 99.505 ;
        RECT 61.320 95.525 62.220 96.425 ;
        RECT 45.835 82.305 46.735 83.205 ;
        RECT 45.860 79.390 46.760 80.290 ;
        RECT 43.500 76.380 44.400 77.280 ;
        RECT 54.820 92.495 55.720 93.395 ;
        RECT 54.845 88.815 55.745 89.715 ;
        RECT 71.345 95.525 72.245 96.425 ;
        RECT 78.510 99.070 79.410 99.970 ;
        RECT 122.020 98.400 122.600 98.980 ;
        RECT 65.315 92.450 66.215 93.350 ;
        RECT 65.080 88.940 65.980 89.840 ;
        RECT 61.320 85.505 62.220 86.405 ;
        RECT 54.820 82.480 55.720 83.380 ;
        RECT 79.235 92.640 80.135 93.540 ;
        RECT 78.510 89.240 79.410 90.140 ;
        RECT 71.345 85.665 72.245 86.565 ;
        RECT 65.315 82.595 66.215 83.495 ;
        RECT 54.845 79.380 55.745 80.280 ;
        RECT 65.080 79.425 65.980 80.325 ;
        RECT 52.350 76.495 52.930 77.075 ;
        RECT 61.320 76.570 62.220 77.470 ;
        RECT 71.345 76.340 72.245 77.240 ;
        RECT 74.360 82.745 75.260 83.645 ;
        RECT 79.200 82.285 80.100 83.185 ;
        RECT 78.670 79.115 79.570 80.015 ;
        RECT 96.505 95.670 97.405 96.570 ;
        RECT 97.960 95.475 98.860 96.375 ;
        RECT 114.835 95.670 115.735 96.570 ;
        RECT 116.290 95.475 117.190 96.375 ;
        RECT 94.600 93.945 95.500 94.845 ;
        RECT 96.030 94.225 96.930 95.125 ;
        RECT 93.570 92.380 94.470 93.280 ;
        RECT 94.980 92.555 95.880 93.455 ;
        RECT 104.635 93.260 105.535 94.160 ;
        RECT 112.930 93.945 113.830 94.845 ;
        RECT 114.360 94.225 115.260 95.125 ;
        RECT 111.900 92.380 112.800 93.280 ;
        RECT 113.310 92.555 114.210 93.455 ;
        RECT 89.665 90.160 90.565 91.060 ;
        RECT 91.220 90.875 92.120 91.775 ;
        RECT 92.865 90.975 93.765 91.875 ;
        RECT 107.995 90.160 108.895 91.060 ;
        RECT 109.550 90.875 110.450 91.775 ;
        RECT 111.195 90.975 112.095 91.875 ;
        RECT 88.005 88.715 88.905 89.615 ;
        RECT 106.335 88.735 107.235 89.635 ;
        RECT 89.665 87.800 90.565 88.700 ;
        RECT 107.995 87.800 108.895 88.700 ;
        RECT 90.540 86.335 91.440 87.235 ;
        RECT 92.000 86.335 92.900 87.235 ;
        RECT 108.870 86.335 109.770 87.235 ;
        RECT 110.330 86.335 111.230 87.235 ;
        RECT 92.615 84.910 93.515 85.810 ;
        RECT 94.105 84.815 95.005 85.715 ;
        RECT 110.945 84.910 111.845 85.810 ;
        RECT 112.435 84.815 113.335 85.715 ;
        RECT 92.615 82.965 93.515 83.865 ;
        RECT 94.310 82.990 95.210 83.890 ;
        RECT 110.945 82.965 111.845 83.865 ;
        RECT 112.640 82.990 113.540 83.890 ;
        RECT 94.885 81.425 95.785 82.325 ;
        RECT 96.390 81.530 97.290 82.430 ;
        RECT 98.040 81.425 98.940 82.325 ;
        RECT 113.215 81.425 114.115 82.325 ;
        RECT 114.720 81.530 115.620 82.430 ;
        RECT 116.370 81.425 117.270 82.325 ;
        RECT 96.265 77.380 97.165 78.280 ;
        RECT 97.670 77.185 98.570 78.085 ;
        RECT 45.835 73.300 46.735 74.200 ;
        RECT 54.820 73.275 55.720 74.175 ;
        RECT 65.315 73.420 66.215 74.320 ;
        RECT 73.955 73.120 74.855 74.020 ;
        RECT 79.330 72.765 80.230 73.665 ;
        RECT 51.545 71.385 52.445 72.285 ;
        RECT 58.270 69.600 58.850 70.180 ;
        RECT 63.540 68.415 64.440 69.315 ;
        RECT 74.360 69.040 74.940 69.620 ;
        RECT 51.430 66.100 52.330 67.000 ;
        RECT 51.545 64.845 52.445 65.745 ;
        RECT 63.540 66.595 64.440 67.495 ;
        RECT 63.540 64.775 64.440 65.675 ;
        RECT 63.550 62.960 64.450 63.860 ;
        RECT 37.410 57.720 37.990 58.300 ;
        RECT 37.410 47.030 37.990 47.610 ;
        RECT 43.635 44.920 44.535 45.820 ;
        RECT 47.830 59.565 48.410 60.145 ;
        RECT 51.430 59.410 52.330 60.310 ;
        RECT 51.545 58.150 52.445 59.050 ;
        RECT 63.550 61.135 64.450 62.035 ;
        RECT 63.550 59.310 64.450 60.210 ;
        RECT 63.540 57.500 64.440 58.400 ;
        RECT 61.245 55.675 62.145 56.575 ;
        RECT 63.550 55.675 64.450 56.575 ;
        RECT 73.040 55.615 73.620 56.195 ;
        RECT 114.865 77.135 115.765 78.035 ;
        RECT 116.320 76.940 117.220 77.840 ;
        RECT 94.310 75.655 95.210 76.555 ;
        RECT 95.740 75.935 96.640 76.835 ;
        RECT 112.960 75.410 113.860 76.310 ;
        RECT 114.390 75.690 115.290 76.590 ;
        RECT 93.280 74.090 94.180 74.990 ;
        RECT 94.690 74.265 95.590 75.165 ;
        RECT 111.930 73.845 112.830 74.745 ;
        RECT 113.340 74.020 114.240 74.920 ;
        RECT 89.375 71.870 90.275 72.770 ;
        RECT 90.930 72.585 91.830 73.485 ;
        RECT 92.575 72.685 93.475 73.585 ;
        RECT 108.025 71.625 108.925 72.525 ;
        RECT 109.580 72.340 110.480 73.240 ;
        RECT 111.225 72.440 112.125 73.340 ;
        RECT 87.715 70.445 88.615 71.345 ;
        RECT 89.375 69.510 90.275 70.410 ;
        RECT 106.365 70.215 107.265 71.115 ;
        RECT 108.025 69.265 108.925 70.165 ;
        RECT 90.250 68.045 91.150 68.945 ;
        RECT 91.710 68.045 92.610 68.945 ;
        RECT 108.900 67.800 109.800 68.700 ;
        RECT 110.360 67.800 111.260 68.700 ;
        RECT 92.325 66.620 93.225 67.520 ;
        RECT 93.815 66.525 94.715 67.425 ;
        RECT 110.975 66.375 111.875 67.275 ;
        RECT 112.465 66.280 113.365 67.180 ;
        RECT 92.325 64.675 93.225 65.575 ;
        RECT 94.020 64.700 94.920 65.600 ;
        RECT 94.595 63.135 95.495 64.035 ;
        RECT 96.100 63.240 97.000 64.140 ;
        RECT 97.750 63.135 98.650 64.035 ;
        RECT 110.975 64.430 111.875 65.330 ;
        RECT 112.670 64.455 113.570 65.355 ;
        RECT 113.245 62.890 114.145 63.790 ;
        RECT 114.750 62.995 115.650 63.895 ;
        RECT 116.400 62.890 117.300 63.790 ;
        RECT 51.430 52.745 52.330 53.645 ;
        RECT 51.470 51.220 52.370 52.120 ;
        RECT 107.015 57.365 107.915 58.265 ;
        RECT 108.600 57.255 109.500 58.155 ;
        RECT 110.020 57.365 110.920 58.265 ;
        RECT 111.600 57.255 112.500 58.155 ;
        RECT 113.990 57.365 114.890 58.265 ;
        RECT 106.350 55.845 107.250 56.745 ;
        RECT 106.015 54.170 106.915 55.070 ;
        RECT 107.570 54.290 108.470 55.190 ;
        RECT 61.445 50.855 62.345 51.755 ;
        RECT 63.775 51.710 64.675 52.610 ;
        RECT 73.040 51.865 73.620 52.445 ;
        RECT 106.530 52.115 107.430 53.015 ;
        RECT 60.090 49.690 60.670 50.270 ;
        RECT 61.445 48.970 62.345 49.870 ;
        RECT 63.775 49.890 64.675 50.790 ;
        RECT 72.980 49.970 73.880 50.870 ;
        RECT 106.015 50.550 106.915 51.450 ;
        RECT 61.445 47.145 62.345 48.045 ;
        RECT 63.775 48.070 64.675 48.970 ;
        RECT 106.530 48.835 107.430 49.735 ;
        RECT 72.920 47.400 73.820 48.300 ;
        RECT 51.430 46.120 52.330 47.020 ;
        RECT 63.785 46.250 64.685 47.150 ;
        RECT 106.015 46.800 106.915 47.700 ;
        RECT 107.570 46.795 108.470 47.695 ;
        RECT 48.210 44.915 49.110 45.815 ;
        RECT 61.445 45.270 62.345 46.170 ;
        RECT 63.785 44.430 64.685 45.330 ;
        RECT 73.030 44.895 73.930 45.795 ;
        RECT 46.710 42.775 47.610 43.675 ;
        RECT 61.445 43.450 62.345 44.350 ;
        RECT 106.690 45.195 107.590 46.095 ;
        RECT 39.355 39.890 40.255 40.790 ;
        RECT 43.655 38.260 44.555 39.160 ;
        RECT 48.165 39.900 49.065 40.800 ;
        RECT 48.210 38.285 49.110 39.185 ;
        RECT 61.445 41.710 62.345 42.610 ;
        RECT 63.785 42.605 64.685 43.505 ;
        RECT 73.030 42.285 73.930 43.185 ;
        RECT 107.570 43.665 108.470 44.565 ;
        RECT 109.100 43.705 110.000 44.605 ;
        RECT 110.470 43.640 111.370 44.540 ;
        RECT 111.830 43.745 112.730 44.645 ;
        RECT 113.990 43.895 114.890 44.795 ;
        RECT 125.330 43.985 125.910 44.565 ;
        RECT 61.445 39.875 62.345 40.775 ;
        RECT 63.775 40.795 64.675 41.695 ;
        RECT 97.225 41.185 98.125 42.085 ;
        RECT 63.785 38.970 64.685 39.870 ;
        RECT 73.030 39.800 73.930 40.700 ;
        RECT 39.005 33.185 39.905 34.085 ;
        RECT 43.615 32.145 44.515 33.045 ;
        RECT 46.710 35.810 47.610 36.710 ;
        RECT 57.670 36.220 58.570 37.120 ;
        RECT 48.150 33.195 49.050 34.095 ;
        RECT 49.400 32.125 50.300 33.025 ;
        RECT 59.005 35.665 59.905 36.565 ;
        RECT 59.005 32.620 59.905 33.520 ;
        RECT 39.005 27.070 39.905 27.970 ;
        RECT 43.655 25.720 44.555 26.620 ;
        RECT 46.710 29.525 47.610 30.425 ;
        RECT 48.185 27.100 49.085 28.000 ;
        RECT 49.400 25.720 50.300 26.620 ;
        RECT 46.710 23.450 47.610 24.350 ;
        RECT 38.015 20.675 38.915 21.575 ;
        RECT 48.140 20.695 49.040 21.595 ;
        RECT 73.075 38.275 73.655 38.855 ;
        RECT 72.845 36.025 73.745 36.925 ;
        RECT 74.305 36.895 74.885 37.475 ;
        RECT 70.750 34.305 71.650 35.205 ;
        RECT 112.660 40.165 113.240 40.745 ;
        RECT 97.225 18.825 98.125 19.725 ;
        RECT 154.730 8.945 155.630 9.845 ;
        RECT 134.415 7.465 135.315 8.365 ;
        RECT 112.305 5.375 113.205 6.275 ;
      LAYER met2 ;
        RECT 56.925 219.620 58.095 219.635 ;
        RECT 56.915 218.620 60.870 219.620 ;
        RECT 56.925 218.505 58.095 218.620 ;
        RECT 132.085 215.935 133.255 215.980 ;
        RECT 127.550 214.935 133.255 215.935 ;
        RECT 132.085 214.850 133.255 214.935 ;
        RECT 7.785 214.705 8.955 214.720 ;
        RECT 7.775 213.705 11.730 214.705 ;
        RECT 7.785 213.590 8.955 213.705 ;
        RECT 97.295 210.005 98.025 210.775 ;
        RECT 105.490 210.145 106.220 210.915 ;
        RECT 102.795 207.445 103.375 207.545 ;
        RECT 106.715 207.445 107.295 207.545 ;
        RECT 63.845 207.165 64.425 207.335 ;
        RECT 92.930 207.165 93.510 207.335 ;
        RECT 102.795 207.305 107.295 207.445 ;
        RECT 63.845 206.865 95.040 207.165 ;
        RECT 102.795 206.905 103.375 207.305 ;
        RECT 63.845 206.695 64.425 206.865 ;
        RECT 92.930 206.695 93.510 206.865 ;
        RECT 53.270 206.205 53.850 206.405 ;
        RECT 53.270 205.905 60.575 206.205 ;
        RECT 53.270 205.765 53.850 205.905 ;
        RECT 53.230 201.365 53.810 201.595 ;
        RECT 60.275 201.365 60.575 205.905 ;
        RECT 63.665 203.380 64.245 203.530 ;
        RECT 92.930 203.380 93.510 203.550 ;
        RECT 63.665 203.080 93.510 203.380 ;
        RECT 63.665 202.890 64.245 203.080 ;
        RECT 92.930 202.910 93.510 203.080 ;
        RECT 63.805 202.415 64.105 202.890 ;
        RECT 63.665 201.775 64.245 202.415 ;
        RECT 53.230 201.065 76.380 201.365 ;
        RECT 53.230 200.955 53.810 201.065 ;
        RECT 76.080 198.125 76.380 201.065 ;
        RECT 75.980 197.485 76.560 198.125 ;
        RECT 52.940 186.525 54.070 187.695 ;
        RECT 56.390 183.640 56.970 184.280 ;
        RECT 54.205 181.760 54.785 181.930 ;
        RECT 56.535 181.760 56.835 183.640 ;
        RECT 54.205 181.460 56.835 181.760 ;
        RECT 54.205 181.290 54.785 181.460 ;
        RECT 88.995 173.150 89.575 173.320 ;
        RECT 88.995 173.110 93.295 173.150 ;
        RECT 94.740 173.110 95.040 206.865 ;
        RECT 97.295 202.830 98.025 203.600 ;
        RECT 102.880 200.230 103.460 200.480 ;
        RECT 105.025 200.230 105.165 207.305 ;
        RECT 106.715 206.905 107.295 207.305 ;
        RECT 105.490 203.065 106.220 203.835 ;
        RECT 106.800 200.230 107.380 200.480 ;
        RECT 102.880 200.090 107.380 200.230 ;
        RECT 102.880 199.840 103.460 200.090 ;
        RECT 97.295 195.880 98.025 196.650 ;
        RECT 102.880 193.350 103.460 193.600 ;
        RECT 105.025 193.350 105.165 200.090 ;
        RECT 106.800 199.840 107.380 200.090 ;
        RECT 105.490 196.195 106.220 196.965 ;
        RECT 106.800 193.350 107.380 193.600 ;
        RECT 102.880 193.210 107.380 193.350 ;
        RECT 102.880 192.960 103.460 193.210 ;
        RECT 95.525 188.805 96.255 189.575 ;
        RECT 97.295 188.855 98.025 189.625 ;
        RECT 97.295 186.190 98.025 186.595 ;
        RECT 102.880 186.190 103.460 186.440 ;
        RECT 105.025 186.190 105.165 193.210 ;
        RECT 106.800 192.960 107.380 193.210 ;
        RECT 105.490 188.855 106.220 189.625 ;
        RECT 106.800 186.190 107.380 186.440 ;
        RECT 97.295 186.050 107.380 186.190 ;
        RECT 97.295 185.825 98.025 186.050 ;
        RECT 102.880 185.800 103.460 186.050 ;
        RECT 106.800 185.800 107.380 186.050 ;
        RECT 88.995 172.850 95.040 173.110 ;
        RECT 88.995 172.680 89.575 172.850 ;
        RECT 92.995 172.810 95.040 172.850 ;
        RECT 89.020 169.135 89.600 169.350 ;
        RECT 85.980 168.835 89.600 169.135 ;
        RECT 52.505 167.260 53.205 167.265 ;
        RECT 52.275 166.560 54.995 167.260 ;
        RECT 52.295 162.580 52.875 162.585 ;
        RECT 54.295 162.580 54.995 166.560 ;
        RECT 52.295 161.945 54.995 162.580 ;
        RECT 52.335 161.880 54.995 161.945 ;
        RECT 52.300 157.820 53.195 157.835 ;
        RECT 54.295 157.820 54.995 161.880 ;
        RECT 85.980 159.205 86.280 168.835 ;
        RECT 89.020 168.710 89.600 168.835 ;
        RECT 89.010 163.090 89.590 163.260 ;
        RECT 92.995 163.090 93.295 172.810 ;
        RECT 105.460 169.790 106.190 170.560 ;
        RECT 93.735 163.090 94.315 163.290 ;
        RECT 89.010 162.790 94.315 163.090 ;
        RECT 105.460 163.000 106.190 163.770 ;
        RECT 89.010 162.620 89.590 162.790 ;
        RECT 93.735 162.650 94.315 162.790 ;
        RECT 85.875 159.190 86.455 159.205 ;
        RECT 89.020 159.190 89.600 159.360 ;
        RECT 85.875 158.890 89.600 159.190 ;
        RECT 85.875 158.565 86.455 158.890 ;
        RECT 89.020 158.720 89.600 158.890 ;
        RECT 55.175 157.820 55.875 157.835 ;
        RECT 52.240 157.120 55.875 157.820 ;
        RECT 111.285 123.655 112.455 123.715 ;
        RECT 111.285 122.655 115.545 123.655 ;
        RECT 111.285 122.585 112.455 122.655 ;
        RECT 7.785 110.795 8.955 110.810 ;
        RECT 7.775 109.795 11.730 110.795 ;
        RECT 137.740 110.345 138.910 110.390 ;
        RECT 53.965 110.190 82.825 110.330 ;
        RECT 7.785 109.680 8.955 109.795 ;
        RECT 45.860 109.275 46.760 109.465 ;
        RECT 43.405 108.575 46.760 109.275 ;
        RECT 43.405 106.950 44.105 108.575 ;
        RECT 45.860 108.505 46.760 108.575 ;
        RECT 53.965 109.065 54.105 110.190 ;
        RECT 54.845 109.065 55.745 109.475 ;
        RECT 53.965 108.925 55.745 109.065 ;
        RECT 43.405 105.990 45.005 106.950 ;
        RECT 43.405 100.600 44.105 105.990 ;
        RECT 45.720 102.235 46.850 103.405 ;
        RECT 45.860 100.600 46.760 100.615 ;
        RECT 43.405 99.900 46.760 100.600 ;
        RECT 43.405 97.155 44.105 99.900 ;
        RECT 45.730 99.865 46.760 99.900 ;
        RECT 45.860 99.655 46.760 99.865 ;
        RECT 53.965 99.015 54.105 108.925 ;
        RECT 54.845 108.515 55.745 108.925 ;
        RECT 64.150 109.065 64.290 110.190 ;
        RECT 65.080 109.065 65.980 109.475 ;
        RECT 73.410 109.225 74.140 109.995 ;
        RECT 78.585 109.940 79.485 110.000 ;
        RECT 78.585 109.240 81.540 109.940 ;
        RECT 64.150 108.925 65.980 109.065 ;
        RECT 78.585 109.040 79.485 109.240 ;
        RECT 61.320 106.675 62.220 106.805 ;
        RECT 61.300 105.845 62.220 106.675 ;
        RECT 54.705 102.270 55.835 103.440 ;
        RECT 54.845 99.015 55.745 99.515 ;
        RECT 53.955 98.875 55.745 99.015 ;
        RECT 43.405 96.195 45.005 97.155 ;
        RECT 37.185 89.580 37.765 89.590 ;
        RECT 43.405 89.580 44.105 96.195 ;
        RECT 45.720 92.325 46.850 93.495 ;
        RECT 37.185 89.395 46.310 89.580 ;
        RECT 37.185 88.950 46.760 89.395 ;
        RECT 53.965 89.335 54.105 98.875 ;
        RECT 54.845 98.555 55.745 98.875 ;
        RECT 61.300 96.455 62.000 105.845 ;
        RECT 64.150 99.035 64.290 108.925 ;
        RECT 65.080 108.515 65.980 108.925 ;
        RECT 80.840 107.985 81.540 109.240 ;
        RECT 80.840 107.285 82.410 107.985 ;
        RECT 71.345 105.845 72.245 106.805 ;
        RECT 65.200 102.210 66.330 103.380 ;
        RECT 65.080 99.035 65.980 99.535 ;
        RECT 64.150 98.895 65.980 99.035 ;
        RECT 61.300 95.495 62.220 96.455 ;
        RECT 54.705 92.360 55.835 93.530 ;
        RECT 54.845 89.335 55.745 89.745 ;
        RECT 53.955 89.195 55.745 89.335 ;
        RECT 37.475 88.880 46.760 88.950 ;
        RECT 43.405 87.795 44.105 88.880 ;
        RECT 45.860 88.435 46.760 88.880 ;
        RECT 43.405 86.835 45.005 87.795 ;
        RECT 43.405 80.150 44.105 86.835 ;
        RECT 45.720 82.170 46.850 83.340 ;
        RECT 45.860 80.150 46.760 80.320 ;
        RECT 43.405 79.450 46.760 80.150 ;
        RECT 53.965 79.870 54.105 89.195 ;
        RECT 54.845 88.785 55.745 89.195 ;
        RECT 61.300 86.435 62.000 95.495 ;
        RECT 64.150 89.460 64.290 98.895 ;
        RECT 65.080 98.575 65.980 98.895 ;
        RECT 71.445 96.455 72.145 105.845 ;
        RECT 79.235 102.960 80.135 103.090 ;
        RECT 79.220 102.130 80.135 102.960 ;
        RECT 79.220 101.990 79.920 102.130 ;
        RECT 80.840 101.990 81.540 107.285 ;
        RECT 81.710 107.270 82.410 107.285 ;
        RECT 82.685 106.215 82.825 110.190 ;
        RECT 133.205 109.345 138.910 110.345 ;
        RECT 137.740 109.260 138.910 109.345 ;
        RECT 82.175 105.825 82.825 106.215 ;
        RECT 82.175 105.575 82.755 105.825 ;
        RECT 78.580 101.290 81.540 101.990 ;
        RECT 78.580 100.000 79.280 101.290 ;
        RECT 78.510 99.040 79.410 100.000 ;
        RECT 71.345 95.495 72.245 96.455 ;
        RECT 65.200 92.315 66.330 93.485 ;
        RECT 65.080 89.460 65.980 89.870 ;
        RECT 64.150 89.320 65.980 89.460 ;
        RECT 61.300 85.475 62.220 86.435 ;
        RECT 54.705 82.345 55.835 83.515 ;
        RECT 54.845 79.870 55.745 80.310 ;
        RECT 53.965 79.730 55.745 79.870 ;
        RECT 43.405 77.310 44.105 79.450 ;
        RECT 45.860 79.360 46.760 79.450 ;
        RECT 54.845 79.350 55.745 79.730 ;
        RECT 61.300 77.500 62.000 85.475 ;
        RECT 64.150 79.900 64.290 89.320 ;
        RECT 65.080 88.910 65.980 89.320 ;
        RECT 71.445 86.595 72.145 95.495 ;
        RECT 79.235 92.610 80.135 93.570 ;
        RECT 79.335 91.715 80.035 92.610 ;
        RECT 80.840 91.715 81.540 101.290 ;
        RECT 121.945 98.305 122.675 99.075 ;
        RECT 95.935 97.165 116.790 97.305 ;
        RECT 95.935 95.155 96.075 97.165 ;
        RECT 96.390 95.535 97.520 96.705 ;
        RECT 98.280 96.405 98.420 97.165 ;
        RECT 97.960 95.445 98.860 96.405 ;
        RECT 94.485 93.810 95.615 94.980 ;
        RECT 95.935 94.605 96.930 95.155 ;
        RECT 96.030 94.195 96.930 94.605 ;
        RECT 78.555 91.015 81.540 91.715 ;
        RECT 90.045 92.590 92.960 92.730 ;
        RECT 90.045 91.090 90.185 92.590 ;
        RECT 78.555 90.170 79.255 91.015 ;
        RECT 78.510 89.210 79.410 90.170 ;
        RECT 71.345 85.635 72.245 86.595 ;
        RECT 65.200 82.460 66.330 83.630 ;
        RECT 65.080 79.900 65.980 80.355 ;
        RECT 64.150 79.760 65.980 79.900 ;
        RECT 65.080 79.395 65.980 79.760 ;
        RECT 43.405 76.480 44.400 77.310 ;
        RECT 43.500 76.350 44.400 76.480 ;
        RECT 52.275 76.400 53.005 77.170 ;
        RECT 61.300 76.540 62.220 77.500 ;
        RECT 71.445 77.270 72.145 85.635 ;
        RECT 74.245 82.610 75.375 83.780 ;
        RECT 79.200 82.255 80.100 83.215 ;
        RECT 79.375 81.520 80.075 82.255 ;
        RECT 80.840 81.520 81.540 91.015 ;
        RECT 89.665 90.130 90.565 91.090 ;
        RECT 91.105 90.740 92.235 91.910 ;
        RECT 92.820 91.905 92.960 92.590 ;
        RECT 93.455 92.245 94.585 93.415 ;
        RECT 94.980 93.075 95.880 93.485 ;
        RECT 96.320 93.075 96.460 94.195 ;
        RECT 94.980 92.935 96.460 93.075 ;
        RECT 94.980 92.525 95.880 92.935 ;
        RECT 92.820 91.690 93.765 91.905 ;
        RECT 95.360 91.690 95.500 92.525 ;
        RECT 92.820 91.550 95.500 91.690 ;
        RECT 92.820 91.355 93.765 91.550 ;
        RECT 92.865 90.945 93.765 91.355 ;
        RECT 87.890 88.580 89.020 89.750 ;
        RECT 90.045 88.730 90.185 90.130 ;
        RECT 89.665 88.320 90.565 88.730 ;
        RECT 89.625 87.770 90.565 88.320 ;
        RECT 89.625 85.540 89.765 87.770 ;
        RECT 90.425 86.200 91.555 87.370 ;
        RECT 92.000 86.820 92.900 87.265 ;
        RECT 92.000 86.680 94.625 86.820 ;
        RECT 92.000 86.305 92.900 86.680 ;
        RECT 92.145 85.540 92.285 86.305 ;
        RECT 89.625 85.400 92.285 85.540 ;
        RECT 91.640 82.260 91.780 85.400 ;
        RECT 92.500 84.775 93.630 85.945 ;
        RECT 94.485 85.745 94.625 86.680 ;
        RECT 94.105 84.785 95.005 85.745 ;
        RECT 92.500 82.830 93.630 84.000 ;
        RECT 94.310 83.510 95.210 83.920 ;
        RECT 94.225 82.960 95.210 83.510 ;
        RECT 94.225 82.260 94.365 82.960 ;
        RECT 91.640 82.120 94.365 82.260 ;
        RECT 78.740 80.820 81.540 81.520 ;
        RECT 78.740 80.045 79.440 80.820 ;
        RECT 78.670 79.085 79.570 80.045 ;
        RECT 45.720 73.165 46.850 74.335 ;
        RECT 54.705 73.140 55.835 74.310 ;
        RECT 51.545 72.295 52.445 72.315 ;
        RECT 50.815 72.155 52.445 72.295 ;
        RECT 50.815 65.730 50.955 72.155 ;
        RECT 51.545 71.355 52.445 72.155 ;
        RECT 61.300 71.305 62.000 76.540 ;
        RECT 71.345 76.310 72.245 77.270 ;
        RECT 65.200 73.285 66.330 74.455 ;
        RECT 71.445 71.305 72.145 76.310 ;
        RECT 73.840 72.985 74.970 74.155 ;
        RECT 79.330 72.735 80.230 73.695 ;
        RECT 79.495 71.305 80.195 72.735 ;
        RECT 80.840 71.305 81.540 80.820 ;
        RECT 93.290 80.520 93.430 82.120 ;
        RECT 94.770 81.290 95.900 82.460 ;
        RECT 96.390 81.500 97.290 82.460 ;
        RECT 96.770 80.520 96.910 81.500 ;
        RECT 97.925 81.290 99.055 82.460 ;
        RECT 93.290 80.380 96.910 80.520 ;
        RECT 104.035 78.770 104.175 97.165 ;
        RECT 114.265 95.155 114.405 97.165 ;
        RECT 114.720 95.535 115.850 96.705 ;
        RECT 116.650 96.405 116.790 97.165 ;
        RECT 116.290 95.445 117.190 96.405 ;
        RECT 104.520 93.125 105.650 94.295 ;
        RECT 112.815 93.810 113.945 94.980 ;
        RECT 114.265 94.605 115.260 95.155 ;
        RECT 114.360 94.195 115.260 94.605 ;
        RECT 108.375 92.590 111.290 92.730 ;
        RECT 108.375 91.090 108.515 92.590 ;
        RECT 107.995 90.130 108.895 91.090 ;
        RECT 109.435 90.740 110.565 91.910 ;
        RECT 111.150 91.905 111.290 92.590 ;
        RECT 111.785 92.245 112.915 93.415 ;
        RECT 113.310 93.075 114.210 93.485 ;
        RECT 114.650 93.075 114.790 94.195 ;
        RECT 113.310 92.935 114.790 93.075 ;
        RECT 113.310 92.525 114.210 92.935 ;
        RECT 111.150 91.690 112.095 91.905 ;
        RECT 113.690 91.690 113.830 92.525 ;
        RECT 111.150 91.550 113.830 91.690 ;
        RECT 111.150 91.355 112.095 91.550 ;
        RECT 111.195 90.945 112.095 91.355 ;
        RECT 106.220 88.600 107.350 89.770 ;
        RECT 108.375 88.730 108.515 90.130 ;
        RECT 107.995 88.320 108.895 88.730 ;
        RECT 107.955 87.770 108.895 88.320 ;
        RECT 107.955 85.540 108.095 87.770 ;
        RECT 108.755 86.200 109.885 87.370 ;
        RECT 110.330 86.820 111.230 87.265 ;
        RECT 110.330 86.680 112.955 86.820 ;
        RECT 110.330 86.305 111.230 86.680 ;
        RECT 110.475 85.540 110.615 86.305 ;
        RECT 107.955 85.400 110.615 85.540 ;
        RECT 109.970 82.260 110.110 85.400 ;
        RECT 110.830 84.775 111.960 85.945 ;
        RECT 112.815 85.745 112.955 86.680 ;
        RECT 112.435 84.785 113.335 85.745 ;
        RECT 110.830 82.830 111.960 84.000 ;
        RECT 112.640 83.510 113.540 83.920 ;
        RECT 112.555 82.960 113.540 83.510 ;
        RECT 112.555 82.260 112.695 82.960 ;
        RECT 109.970 82.120 112.695 82.260 ;
        RECT 111.620 80.520 111.760 82.120 ;
        RECT 113.100 81.290 114.230 82.460 ;
        RECT 114.720 81.500 115.620 82.460 ;
        RECT 115.100 80.520 115.240 81.500 ;
        RECT 116.255 81.290 117.385 82.460 ;
        RECT 111.620 80.380 115.240 80.520 ;
        RECT 95.860 78.630 116.780 78.770 ;
        RECT 95.860 76.865 96.000 78.630 ;
        RECT 96.150 77.245 97.280 78.415 ;
        RECT 97.875 78.115 98.015 78.630 ;
        RECT 97.670 77.155 98.570 78.115 ;
        RECT 94.195 75.520 95.325 76.690 ;
        RECT 95.740 75.905 96.640 76.865 ;
        RECT 114.295 76.620 114.435 78.630 ;
        RECT 114.750 77.000 115.880 78.170 ;
        RECT 116.640 77.870 116.780 78.630 ;
        RECT 116.320 76.910 117.220 77.870 ;
        RECT 89.755 74.300 92.670 74.440 ;
        RECT 89.755 72.800 89.895 74.300 ;
        RECT 89.375 71.840 90.275 72.800 ;
        RECT 90.815 72.450 91.945 73.620 ;
        RECT 92.530 73.615 92.670 74.300 ;
        RECT 93.165 73.955 94.295 75.125 ;
        RECT 94.690 74.785 95.590 75.195 ;
        RECT 96.030 74.785 96.170 75.905 ;
        RECT 112.845 75.275 113.975 76.445 ;
        RECT 114.295 76.070 115.290 76.620 ;
        RECT 114.390 75.660 115.290 76.070 ;
        RECT 94.690 74.645 96.170 74.785 ;
        RECT 94.690 74.235 95.590 74.645 ;
        RECT 92.530 73.400 93.475 73.615 ;
        RECT 95.070 73.400 95.210 74.235 ;
        RECT 92.530 73.260 95.210 73.400 ;
        RECT 108.405 74.055 111.320 74.195 ;
        RECT 92.530 73.065 93.475 73.260 ;
        RECT 92.575 72.655 93.475 73.065 ;
        RECT 108.405 72.555 108.545 74.055 ;
        RECT 61.300 70.605 81.540 71.305 ;
        RECT 58.195 69.505 58.925 70.275 ;
        RECT 62.925 68.935 63.065 70.605 ;
        RECT 63.540 68.935 64.440 69.345 ;
        RECT 74.300 69.010 75.000 70.605 ;
        RECT 87.600 70.310 88.730 71.480 ;
        RECT 89.755 70.440 89.895 71.840 ;
        RECT 108.025 71.595 108.925 72.555 ;
        RECT 109.465 72.205 110.595 73.375 ;
        RECT 111.180 73.370 111.320 74.055 ;
        RECT 111.815 73.710 112.945 74.880 ;
        RECT 113.340 74.540 114.240 74.950 ;
        RECT 114.680 74.540 114.820 75.660 ;
        RECT 113.340 74.400 114.820 74.540 ;
        RECT 113.340 73.990 114.240 74.400 ;
        RECT 111.180 73.155 112.125 73.370 ;
        RECT 113.720 73.155 113.860 73.990 ;
        RECT 111.180 73.015 113.860 73.155 ;
        RECT 111.180 72.820 112.125 73.015 ;
        RECT 111.225 72.410 112.125 72.820 ;
        RECT 89.375 70.030 90.275 70.440 ;
        RECT 106.250 70.080 107.380 71.250 ;
        RECT 108.405 70.195 108.545 71.595 ;
        RECT 89.335 69.480 90.275 70.030 ;
        RECT 108.025 69.785 108.925 70.195 ;
        RECT 62.925 68.795 64.440 68.935 ;
        RECT 51.315 65.965 52.445 67.135 ;
        RECT 62.925 66.965 63.065 68.795 ;
        RECT 63.540 68.385 64.440 68.795 ;
        RECT 63.540 66.965 64.440 67.525 ;
        RECT 62.925 66.825 64.440 66.965 ;
        RECT 89.335 66.875 89.475 69.480 ;
        RECT 107.985 69.235 108.925 69.785 ;
        RECT 90.135 67.910 91.265 69.080 ;
        RECT 91.710 68.155 92.610 68.975 ;
        RECT 91.710 68.015 94.335 68.155 ;
        RECT 91.855 66.875 91.995 68.015 ;
        RECT 51.545 65.730 52.445 65.775 ;
        RECT 50.815 65.590 52.445 65.730 ;
        RECT 47.755 59.470 48.485 60.240 ;
        RECT 50.815 59.010 50.955 65.590 ;
        RECT 51.545 64.815 52.445 65.590 ;
        RECT 62.925 65.315 63.065 66.825 ;
        RECT 63.540 66.565 64.440 66.825 ;
        RECT 85.260 66.735 91.995 66.875 ;
        RECT 63.540 65.315 64.440 65.705 ;
        RECT 62.925 65.175 64.440 65.315 ;
        RECT 62.925 63.450 63.065 65.175 ;
        RECT 63.540 64.745 64.440 65.175 ;
        RECT 63.550 63.450 64.450 63.890 ;
        RECT 62.925 63.310 64.450 63.450 ;
        RECT 62.925 61.645 63.065 63.310 ;
        RECT 63.550 62.930 64.450 63.310 ;
        RECT 63.550 61.645 64.450 62.065 ;
        RECT 62.925 61.505 64.450 61.645 ;
        RECT 51.315 59.275 52.445 60.445 ;
        RECT 62.925 59.820 63.065 61.505 ;
        RECT 63.550 61.105 64.450 61.505 ;
        RECT 63.550 59.820 64.450 60.240 ;
        RECT 62.925 59.680 64.450 59.820 ;
        RECT 51.545 59.010 52.445 59.080 ;
        RECT 50.815 58.870 52.445 59.010 ;
        RECT 50.815 58.360 50.955 58.870 ;
        RECT 37.410 57.660 50.955 58.360 ;
        RECT 51.545 58.120 52.445 58.870 ;
        RECT 50.815 52.120 50.955 57.660 ;
        RECT 62.925 57.895 63.065 59.680 ;
        RECT 63.550 59.280 64.450 59.680 ;
        RECT 63.540 57.895 64.440 58.430 ;
        RECT 62.925 57.755 64.440 57.895 ;
        RECT 61.245 55.645 62.145 56.605 ;
        RECT 62.925 56.270 63.065 57.755 ;
        RECT 63.540 57.470 64.440 57.755 ;
        RECT 63.550 56.270 64.450 56.605 ;
        RECT 62.925 56.130 64.450 56.270 ;
        RECT 63.550 55.645 64.450 56.130 ;
        RECT 61.625 54.135 61.765 55.645 ;
        RECT 72.965 55.520 73.695 56.290 ;
        RECT 61.625 53.995 64.275 54.135 ;
        RECT 51.315 52.610 52.445 53.780 ;
        RECT 64.135 52.640 64.275 53.995 ;
        RECT 63.775 52.240 64.675 52.640 ;
        RECT 51.470 52.120 52.370 52.150 ;
        RECT 50.815 51.980 52.370 52.120 ;
        RECT 51.470 51.190 52.370 51.980 ;
        RECT 63.160 52.100 64.675 52.240 ;
        RECT 61.330 50.720 62.460 51.890 ;
        RECT 59.815 49.395 60.945 50.565 ;
        RECT 63.160 50.260 63.300 52.100 ;
        RECT 63.775 51.680 64.675 52.100 ;
        RECT 72.965 51.770 73.695 52.540 ;
        RECT 63.775 50.260 64.675 50.820 ;
        RECT 63.160 50.120 64.675 50.260 ;
        RECT 61.330 48.835 62.460 50.005 ;
        RECT 63.160 48.610 63.300 50.120 ;
        RECT 63.775 49.860 64.675 50.120 ;
        RECT 72.865 49.835 73.995 51.005 ;
        RECT 63.775 48.610 64.675 49.000 ;
        RECT 63.160 48.470 64.675 48.610 ;
        RECT 37.350 47.590 38.050 47.640 ;
        RECT 37.350 46.890 44.435 47.590 ;
        RECT 43.735 45.850 44.435 46.890 ;
        RECT 51.315 45.985 52.445 47.155 ;
        RECT 61.330 47.010 62.460 48.180 ;
        RECT 63.160 46.745 63.300 48.470 ;
        RECT 63.775 48.040 64.675 48.470 ;
        RECT 72.805 47.265 73.935 48.435 ;
        RECT 63.785 46.745 64.685 47.180 ;
        RECT 63.160 46.605 64.685 46.745 ;
        RECT 43.635 45.715 44.535 45.850 ;
        RECT 48.210 45.730 49.110 45.845 ;
        RECT 48.210 45.715 56.665 45.730 ;
        RECT 43.635 45.030 56.665 45.715 ;
        RECT 61.330 45.135 62.460 46.305 ;
        RECT 43.635 45.015 49.110 45.030 ;
        RECT 43.635 44.890 44.535 45.015 ;
        RECT 39.240 39.755 40.370 40.925 ;
        RECT 43.655 38.860 44.555 39.190 ;
        RECT 44.765 38.860 44.905 45.015 ;
        RECT 43.655 38.560 44.905 38.860 ;
        RECT 43.655 38.230 44.555 38.560 ;
        RECT 38.890 33.050 40.020 34.220 ;
        RECT 43.615 32.540 44.515 33.075 ;
        RECT 44.765 32.540 44.905 38.560 ;
        RECT 43.615 32.240 44.905 32.540 ;
        RECT 43.615 32.115 44.515 32.240 ;
        RECT 38.890 26.935 40.020 28.105 ;
        RECT 43.655 26.050 44.555 26.650 ;
        RECT 44.765 26.050 44.905 32.240 ;
        RECT 43.655 25.910 44.905 26.050 ;
        RECT 46.210 43.375 46.510 45.015 ;
        RECT 48.210 44.885 49.110 45.015 ;
        RECT 46.710 43.375 47.610 43.705 ;
        RECT 46.210 43.075 47.610 43.375 ;
        RECT 46.210 38.885 46.510 43.075 ;
        RECT 46.710 42.745 47.610 43.075 ;
        RECT 48.050 39.765 49.180 40.935 ;
        RECT 48.210 38.885 49.110 39.215 ;
        RECT 46.210 38.585 49.110 38.885 ;
        RECT 46.210 36.410 46.510 38.585 ;
        RECT 48.210 38.255 49.110 38.585 ;
        RECT 55.965 37.020 56.665 45.030 ;
        RECT 63.160 44.940 63.300 46.605 ;
        RECT 63.785 46.220 64.685 46.605 ;
        RECT 63.785 44.940 64.685 45.360 ;
        RECT 63.160 44.800 64.685 44.940 ;
        RECT 61.330 43.315 62.460 44.485 ;
        RECT 63.160 43.115 63.300 44.800 ;
        RECT 63.785 44.400 64.685 44.800 ;
        RECT 72.915 44.760 74.045 45.930 ;
        RECT 63.785 43.115 64.685 43.535 ;
        RECT 63.160 42.975 64.685 43.115 ;
        RECT 61.330 41.575 62.460 42.745 ;
        RECT 63.160 41.310 63.300 42.975 ;
        RECT 63.785 42.575 64.685 42.975 ;
        RECT 72.915 42.150 74.045 43.320 ;
        RECT 63.775 41.310 64.675 41.725 ;
        RECT 63.160 41.170 64.675 41.310 ;
        RECT 61.330 39.740 62.460 40.910 ;
        RECT 63.160 39.490 63.300 41.170 ;
        RECT 63.775 40.765 64.675 41.170 ;
        RECT 63.785 39.490 64.685 39.900 ;
        RECT 72.915 39.665 74.045 40.835 ;
        RECT 63.160 39.350 64.685 39.490 ;
        RECT 63.785 38.940 64.685 39.350 ;
        RECT 73.000 38.180 73.730 38.950 ;
        RECT 85.260 38.430 85.400 66.735 ;
        RECT 91.520 64.020 91.660 66.735 ;
        RECT 92.210 66.485 93.340 67.655 ;
        RECT 94.195 67.455 94.335 68.015 ;
        RECT 93.815 66.495 94.715 67.455 ;
        RECT 107.985 67.005 108.125 69.235 ;
        RECT 108.785 67.665 109.915 68.835 ;
        RECT 110.360 68.285 111.260 68.730 ;
        RECT 110.360 68.145 112.985 68.285 ;
        RECT 110.360 67.770 111.260 68.145 ;
        RECT 110.505 67.005 110.645 67.770 ;
        RECT 107.985 66.865 110.645 67.005 ;
        RECT 92.210 64.540 93.340 65.710 ;
        RECT 94.020 65.220 94.920 65.630 ;
        RECT 93.730 65.080 94.920 65.220 ;
        RECT 93.730 64.020 93.870 65.080 ;
        RECT 94.020 64.670 94.920 65.080 ;
        RECT 91.520 63.880 93.870 64.020 ;
        RECT 93.000 61.855 93.140 63.880 ;
        RECT 94.480 63.000 95.610 64.170 ;
        RECT 96.100 63.210 97.000 64.170 ;
        RECT 96.480 61.855 96.620 63.210 ;
        RECT 97.635 63.000 98.765 64.170 ;
        RECT 110.000 63.725 110.140 66.865 ;
        RECT 110.860 66.240 111.990 67.410 ;
        RECT 112.845 67.210 112.985 68.145 ;
        RECT 112.465 66.250 113.365 67.210 ;
        RECT 110.860 64.295 111.990 65.465 ;
        RECT 112.670 64.975 113.570 65.385 ;
        RECT 112.585 64.425 113.570 64.975 ;
        RECT 112.585 63.725 112.725 64.425 ;
        RECT 110.000 63.585 112.725 63.725 ;
        RECT 93.000 61.715 96.620 61.855 ;
        RECT 111.650 61.985 111.790 63.585 ;
        RECT 113.130 62.755 114.260 63.925 ;
        RECT 114.750 62.965 115.650 63.925 ;
        RECT 115.130 61.985 115.270 62.965 ;
        RECT 116.285 62.755 117.415 63.925 ;
        RECT 111.650 61.845 115.270 61.985 ;
        RECT 96.480 61.620 96.620 61.715 ;
        RECT 96.480 61.480 96.660 61.620 ;
        RECT 96.520 60.565 96.660 61.480 ;
        RECT 96.520 60.425 103.600 60.565 ;
        RECT 97.110 41.050 98.240 42.220 ;
        RECT 103.460 40.525 103.600 60.425 ;
        RECT 107.115 58.825 114.790 59.525 ;
        RECT 107.115 58.295 107.815 58.825 ;
        RECT 110.145 58.295 110.845 58.825 ;
        RECT 114.090 58.295 114.790 58.825 ;
        RECT 107.015 58.165 107.915 58.295 ;
        RECT 104.585 57.465 107.915 58.165 ;
        RECT 104.585 52.915 105.285 57.465 ;
        RECT 107.015 57.335 107.915 57.465 ;
        RECT 108.485 57.120 109.615 58.290 ;
        RECT 110.020 57.335 110.920 58.295 ;
        RECT 111.485 57.120 112.615 58.290 ;
        RECT 113.990 57.335 114.890 58.295 ;
        RECT 106.235 55.710 107.365 56.880 ;
        RECT 105.900 54.035 107.030 55.205 ;
        RECT 107.570 54.260 108.470 55.220 ;
        RECT 107.770 53.240 108.470 54.260 ;
        RECT 106.630 53.045 108.470 53.240 ;
        RECT 106.530 52.915 108.470 53.045 ;
        RECT 104.525 52.540 108.470 52.915 ;
        RECT 104.525 52.215 107.430 52.540 ;
        RECT 104.525 49.635 105.225 52.215 ;
        RECT 106.530 52.085 107.430 52.215 ;
        RECT 105.900 50.415 107.030 51.585 ;
        RECT 106.530 49.635 107.430 49.765 ;
        RECT 104.525 49.430 107.430 49.635 ;
        RECT 104.510 48.935 107.430 49.430 ;
        RECT 104.510 48.730 105.225 48.935 ;
        RECT 106.530 48.805 107.430 48.935 ;
        RECT 104.510 43.105 105.210 48.730 ;
        RECT 105.900 46.665 107.030 47.835 ;
        RECT 107.570 46.765 108.470 47.725 ;
        RECT 106.575 45.060 107.705 46.230 ;
        RECT 107.950 44.595 108.090 46.765 ;
        RECT 107.570 43.635 108.470 44.595 ;
        RECT 107.935 43.105 108.075 43.635 ;
        RECT 108.985 43.570 110.115 44.740 ;
        RECT 110.470 43.610 111.370 44.570 ;
        RECT 111.715 43.610 112.845 44.780 ;
        RECT 113.990 44.645 114.890 44.825 ;
        RECT 113.990 44.595 125.695 44.645 ;
        RECT 113.990 43.955 125.920 44.595 ;
        RECT 113.990 43.945 125.695 43.955 ;
        RECT 113.990 43.865 114.890 43.945 ;
        RECT 104.510 42.860 108.425 43.105 ;
        RECT 110.535 42.860 111.235 43.610 ;
        RECT 114.090 42.860 114.790 43.865 ;
        RECT 104.510 42.405 114.790 42.860 ;
        RECT 108.005 42.160 114.790 42.405 ;
        RECT 112.650 40.525 113.250 40.775 ;
        RECT 103.460 40.385 113.250 40.525 ;
        RECT 112.650 40.135 113.250 40.385 ;
        RECT 85.240 38.290 85.400 38.430 ;
        RECT 57.985 37.430 71.550 38.130 ;
        RECT 57.985 37.150 58.685 37.430 ;
        RECT 57.670 37.020 58.685 37.150 ;
        RECT 46.710 36.410 47.610 36.740 ;
        RECT 46.210 36.110 47.610 36.410 ;
        RECT 55.965 36.320 58.685 37.020 ;
        RECT 57.670 36.190 58.570 36.320 ;
        RECT 46.210 32.365 46.510 36.110 ;
        RECT 46.710 35.780 47.610 36.110 ;
        RECT 58.890 35.530 60.020 36.700 ;
        RECT 70.850 35.235 71.550 37.430 ;
        RECT 74.305 37.310 74.885 37.505 ;
        RECT 85.240 37.310 85.380 38.290 ;
        RECT 74.305 37.170 85.380 37.310 ;
        RECT 72.730 35.890 73.860 37.060 ;
        RECT 74.305 36.865 74.885 37.170 ;
        RECT 70.750 34.275 71.650 35.235 ;
        RECT 48.035 33.060 49.165 34.230 ;
        RECT 49.400 32.365 50.300 33.055 ;
        RECT 58.890 32.485 60.020 33.655 ;
        RECT 46.210 32.225 50.300 32.365 ;
        RECT 46.210 30.125 46.510 32.225 ;
        RECT 49.400 32.095 50.300 32.225 ;
        RECT 46.710 30.125 47.610 30.455 ;
        RECT 46.210 29.825 47.610 30.125 ;
        RECT 46.210 26.255 46.510 29.825 ;
        RECT 46.710 29.495 47.610 29.825 ;
        RECT 48.070 26.965 49.200 28.135 ;
        RECT 49.400 26.255 50.300 26.650 ;
        RECT 46.210 25.955 50.300 26.255 ;
        RECT 43.655 25.690 44.555 25.910 ;
        RECT 47.010 24.380 47.310 25.955 ;
        RECT 49.400 25.690 50.300 25.955 ;
        RECT 46.710 23.420 47.610 24.380 ;
        RECT 37.900 20.540 39.030 21.710 ;
        RECT 48.025 20.560 49.155 21.730 ;
        RECT 97.110 18.690 98.240 19.860 ;
        RECT 112.255 4.210 113.255 6.275 ;
        RECT 134.365 4.550 135.365 8.365 ;
        RECT 112.215 3.080 113.385 4.210 ;
        RECT 134.190 4.025 135.365 4.550 ;
        RECT 154.680 4.550 155.680 9.845 ;
        RECT 134.190 3.420 135.360 4.025 ;
        RECT 154.680 3.855 155.915 4.550 ;
        RECT 154.745 3.420 155.915 3.855 ;
      LAYER via2 ;
        RECT 56.970 218.530 58.050 219.610 ;
        RECT 132.130 214.875 133.210 215.955 ;
        RECT 7.830 213.615 8.910 214.695 ;
        RECT 97.320 210.050 98.000 210.730 ;
        RECT 105.515 210.190 106.195 210.870 ;
        RECT 52.965 186.570 54.045 187.650 ;
        RECT 97.320 202.875 98.000 203.555 ;
        RECT 105.515 203.110 106.195 203.790 ;
        RECT 97.320 195.925 98.000 196.605 ;
        RECT 105.515 196.240 106.195 196.920 ;
        RECT 95.550 188.850 96.230 189.530 ;
        RECT 97.320 188.900 98.000 189.580 ;
        RECT 97.320 185.870 98.000 186.550 ;
        RECT 105.515 188.900 106.195 189.580 ;
        RECT 105.485 169.835 106.165 170.515 ;
        RECT 105.485 163.045 106.165 163.725 ;
        RECT 111.330 122.610 112.410 123.690 ;
        RECT 7.830 109.705 8.910 110.785 ;
        RECT 45.745 102.280 46.825 103.360 ;
        RECT 73.435 109.270 74.115 109.950 ;
        RECT 54.730 102.315 55.810 103.395 ;
        RECT 45.745 92.370 46.825 93.450 ;
        RECT 65.225 102.255 66.305 103.335 ;
        RECT 54.730 92.405 55.810 93.485 ;
        RECT 45.745 82.215 46.825 83.295 ;
        RECT 137.785 109.285 138.865 110.365 ;
        RECT 65.225 92.360 66.305 93.440 ;
        RECT 54.730 82.390 55.810 83.470 ;
        RECT 121.970 98.350 122.650 99.030 ;
        RECT 96.415 95.580 97.495 96.660 ;
        RECT 94.510 93.855 95.590 94.935 ;
        RECT 65.225 82.505 66.305 83.585 ;
        RECT 52.300 76.445 52.980 77.125 ;
        RECT 74.270 82.655 75.350 83.735 ;
        RECT 91.130 90.785 92.210 91.865 ;
        RECT 93.480 92.290 94.560 93.370 ;
        RECT 87.915 88.625 88.995 89.705 ;
        RECT 90.450 86.245 91.530 87.325 ;
        RECT 92.525 84.820 93.605 85.900 ;
        RECT 92.525 82.875 93.605 83.955 ;
        RECT 45.745 73.210 46.825 74.290 ;
        RECT 54.730 73.185 55.810 74.265 ;
        RECT 65.225 73.330 66.305 74.410 ;
        RECT 73.865 73.030 74.945 74.110 ;
        RECT 94.795 81.335 95.875 82.415 ;
        RECT 97.950 81.335 99.030 82.415 ;
        RECT 114.745 95.580 115.825 96.660 ;
        RECT 104.545 93.170 105.625 94.250 ;
        RECT 112.840 93.855 113.920 94.935 ;
        RECT 109.460 90.785 110.540 91.865 ;
        RECT 111.810 92.290 112.890 93.370 ;
        RECT 106.245 88.645 107.325 89.725 ;
        RECT 108.780 86.245 109.860 87.325 ;
        RECT 110.855 84.820 111.935 85.900 ;
        RECT 110.855 82.875 111.935 83.955 ;
        RECT 113.125 81.335 114.205 82.415 ;
        RECT 116.280 81.335 117.360 82.415 ;
        RECT 96.175 77.290 97.255 78.370 ;
        RECT 94.220 75.565 95.300 76.645 ;
        RECT 114.775 77.045 115.855 78.125 ;
        RECT 90.840 72.495 91.920 73.575 ;
        RECT 93.190 74.000 94.270 75.080 ;
        RECT 112.870 75.320 113.950 76.400 ;
        RECT 58.220 69.550 58.900 70.230 ;
        RECT 87.625 70.355 88.705 71.435 ;
        RECT 109.490 72.250 110.570 73.330 ;
        RECT 111.840 73.755 112.920 74.835 ;
        RECT 106.275 70.125 107.355 71.205 ;
        RECT 51.340 66.010 52.420 67.090 ;
        RECT 90.160 67.955 91.240 69.035 ;
        RECT 47.780 59.515 48.460 60.195 ;
        RECT 51.340 59.320 52.420 60.400 ;
        RECT 72.990 55.565 73.670 56.245 ;
        RECT 51.340 52.655 52.420 53.735 ;
        RECT 61.355 50.765 62.435 51.845 ;
        RECT 59.840 49.440 60.920 50.520 ;
        RECT 72.990 51.815 73.670 52.495 ;
        RECT 61.355 48.880 62.435 49.960 ;
        RECT 72.890 49.880 73.970 50.960 ;
        RECT 51.340 46.030 52.420 47.110 ;
        RECT 61.355 47.055 62.435 48.135 ;
        RECT 72.830 47.310 73.910 48.390 ;
        RECT 61.355 45.180 62.435 46.260 ;
        RECT 39.265 39.800 40.345 40.880 ;
        RECT 38.915 33.095 39.995 34.175 ;
        RECT 38.915 26.980 39.995 28.060 ;
        RECT 48.075 39.810 49.155 40.890 ;
        RECT 61.355 43.360 62.435 44.440 ;
        RECT 72.940 44.805 74.020 45.885 ;
        RECT 61.355 41.620 62.435 42.700 ;
        RECT 72.940 42.195 74.020 43.275 ;
        RECT 61.355 39.785 62.435 40.865 ;
        RECT 72.940 39.710 74.020 40.790 ;
        RECT 73.025 38.225 73.705 38.905 ;
        RECT 92.235 66.530 93.315 67.610 ;
        RECT 108.810 67.710 109.890 68.790 ;
        RECT 92.235 64.585 93.315 65.665 ;
        RECT 94.505 63.045 95.585 64.125 ;
        RECT 97.660 63.045 98.740 64.125 ;
        RECT 110.885 66.285 111.965 67.365 ;
        RECT 110.885 64.340 111.965 65.420 ;
        RECT 113.155 62.800 114.235 63.880 ;
        RECT 116.310 62.800 117.390 63.880 ;
        RECT 97.135 41.095 98.215 42.175 ;
        RECT 108.510 57.165 109.590 58.245 ;
        RECT 111.510 57.165 112.590 58.245 ;
        RECT 106.260 55.755 107.340 56.835 ;
        RECT 105.925 54.080 107.005 55.160 ;
        RECT 105.925 50.460 107.005 51.540 ;
        RECT 105.925 46.710 107.005 47.790 ;
        RECT 106.600 45.105 107.680 46.185 ;
        RECT 109.010 43.615 110.090 44.695 ;
        RECT 111.740 43.655 112.820 44.735 ;
        RECT 58.915 35.575 59.995 36.655 ;
        RECT 72.755 35.935 73.835 37.015 ;
        RECT 48.060 33.105 49.140 34.185 ;
        RECT 58.915 32.530 59.995 33.610 ;
        RECT 48.095 27.010 49.175 28.090 ;
        RECT 37.925 20.585 39.005 21.665 ;
        RECT 48.050 20.605 49.130 21.685 ;
        RECT 97.135 18.735 98.215 19.815 ;
        RECT 112.260 3.105 113.340 4.185 ;
        RECT 134.235 3.445 135.315 4.525 ;
        RECT 154.790 3.445 155.870 4.525 ;
      LAYER met3 ;
        RECT 56.925 219.630 58.095 219.635 ;
        RECT 56.920 218.510 58.100 219.630 ;
        RECT 56.925 218.505 58.095 218.510 ;
        RECT 132.085 215.975 133.255 215.980 ;
        RECT 132.080 214.855 133.260 215.975 ;
        RECT 132.085 214.850 133.255 214.855 ;
        RECT 7.785 214.715 8.955 214.720 ;
        RECT 7.780 213.595 8.960 214.715 ;
        RECT 7.785 213.590 8.955 213.595 ;
        RECT 97.510 210.775 97.810 210.780 ;
        RECT 97.295 210.005 98.025 210.775 ;
        RECT 105.490 210.145 106.220 210.915 ;
        RECT 97.510 206.605 97.810 210.005 ;
        RECT 105.705 206.605 106.005 210.145 ;
        RECT 97.510 206.305 106.005 206.605 ;
        RECT 97.510 203.600 97.810 206.305 ;
        RECT 105.705 203.835 106.005 206.305 ;
        RECT 97.295 202.830 98.025 203.600 ;
        RECT 105.490 203.065 106.220 203.835 ;
        RECT 97.510 196.650 97.810 202.830 ;
        RECT 105.705 196.965 106.005 203.065 ;
        RECT 97.295 195.880 98.025 196.650 ;
        RECT 105.490 196.195 106.220 196.965 ;
        RECT 97.510 189.625 97.810 195.880 ;
        RECT 105.705 189.625 106.005 196.195 ;
        RECT 95.525 189.340 96.255 189.575 ;
        RECT 97.295 189.340 98.025 189.625 ;
        RECT 95.525 189.040 98.025 189.340 ;
        RECT 95.525 188.805 96.255 189.040 ;
        RECT 97.295 188.855 98.025 189.040 ;
        RECT 105.490 188.855 106.220 189.625 ;
        RECT 52.940 187.195 54.070 187.695 ;
        RECT 52.940 186.895 57.215 187.195 ;
        RECT 52.940 186.525 54.070 186.895 ;
        RECT 56.915 185.395 57.215 186.895 ;
        RECT 97.295 185.825 98.025 186.595 ;
        RECT 97.510 185.395 97.810 185.825 ;
        RECT 56.915 185.095 97.810 185.395 ;
        RECT 105.705 170.560 106.005 188.855 ;
        RECT 105.460 169.790 106.190 170.560 ;
        RECT 105.705 163.770 106.005 169.790 ;
        RECT 105.460 163.000 106.190 163.770 ;
        RECT 111.285 123.710 112.455 123.715 ;
        RECT 111.280 122.590 112.460 123.710 ;
        RECT 111.285 122.585 112.455 122.590 ;
        RECT 7.785 110.805 8.955 110.810 ;
        RECT 7.780 109.685 8.960 110.805 ;
        RECT 137.740 110.385 138.910 110.390 ;
        RECT 73.410 109.875 74.140 109.995 ;
        RECT 44.050 109.860 74.140 109.875 ;
        RECT 7.785 109.680 8.955 109.685 ;
        RECT 42.700 109.575 74.140 109.860 ;
        RECT 42.700 109.560 44.350 109.575 ;
        RECT 42.700 102.655 43.000 109.560 ;
        RECT 73.410 109.225 74.140 109.575 ;
        RECT 137.735 109.265 138.915 110.385 ;
        RECT 137.740 109.260 138.910 109.265 ;
        RECT 45.720 102.655 46.850 103.405 ;
        RECT 42.700 102.355 46.850 102.655 ;
        RECT 42.700 92.785 43.000 102.355 ;
        RECT 45.720 102.235 46.850 102.355 ;
        RECT 54.705 102.270 55.835 103.440 ;
        RECT 55.120 100.765 55.420 102.270 ;
        RECT 65.200 102.210 66.330 103.380 ;
        RECT 65.385 101.190 65.685 102.210 ;
        RECT 53.455 100.465 55.420 100.765 ;
        RECT 63.820 100.890 65.765 101.190 ;
        RECT 45.720 92.785 46.850 93.495 ;
        RECT 42.700 92.485 46.850 92.785 ;
        RECT 45.720 92.325 46.850 92.485 ;
        RECT 53.455 93.205 53.755 100.465 ;
        RECT 54.705 93.205 55.835 93.530 ;
        RECT 53.455 92.905 55.835 93.205 ;
        RECT 45.720 82.690 46.850 83.340 ;
        RECT 44.755 82.390 46.850 82.690 ;
        RECT 44.755 73.780 45.055 82.390 ;
        RECT 45.720 82.170 46.850 82.390 ;
        RECT 53.455 83.080 53.755 92.905 ;
        RECT 54.705 92.360 55.835 92.905 ;
        RECT 63.820 92.925 64.120 100.890 ;
        RECT 121.945 99.040 122.675 99.075 ;
        RECT 104.695 98.340 122.675 99.040 ;
        RECT 96.390 96.510 97.520 96.705 ;
        RECT 94.700 95.810 97.520 96.510 ;
        RECT 94.700 94.980 95.400 95.810 ;
        RECT 96.390 95.535 97.520 95.810 ;
        RECT 94.485 94.755 95.615 94.980 ;
        RECT 93.365 94.055 95.615 94.755 ;
        RECT 104.695 94.295 105.395 98.340 ;
        RECT 121.945 98.305 122.675 98.340 ;
        RECT 114.720 96.510 115.850 96.705 ;
        RECT 113.030 95.810 115.850 96.510 ;
        RECT 113.030 94.980 113.730 95.810 ;
        RECT 114.720 95.535 115.850 95.810 ;
        RECT 112.815 94.755 113.945 94.980 ;
        RECT 65.200 92.925 66.330 93.485 ;
        RECT 93.365 93.415 94.065 94.055 ;
        RECT 94.485 93.810 95.615 94.055 ;
        RECT 93.365 93.400 94.585 93.415 ;
        RECT 63.820 92.625 66.330 92.925 ;
        RECT 54.705 83.080 55.835 83.515 ;
        RECT 53.455 82.780 55.835 83.080 ;
        RECT 52.275 76.935 53.005 77.170 ;
        RECT 53.455 76.935 53.755 82.780 ;
        RECT 54.705 82.345 55.835 82.780 ;
        RECT 63.820 83.175 64.120 92.625 ;
        RECT 65.200 92.315 66.330 92.625 ;
        RECT 91.320 92.700 94.585 93.400 ;
        RECT 104.520 93.125 105.650 94.295 ;
        RECT 111.780 94.055 113.945 94.755 ;
        RECT 111.780 93.485 112.480 94.055 ;
        RECT 112.815 93.810 113.945 94.055 ;
        RECT 109.650 93.415 112.700 93.485 ;
        RECT 91.320 91.910 92.020 92.700 ;
        RECT 93.455 92.245 94.585 92.700 ;
        RECT 109.650 92.785 112.915 93.415 ;
        RECT 109.650 91.910 110.350 92.785 ;
        RECT 111.785 92.245 112.915 92.785 ;
        RECT 91.105 91.530 92.235 91.910 ;
        RECT 109.435 91.615 110.565 91.910 ;
        RECT 88.150 90.830 92.235 91.530 ;
        RECT 88.150 89.750 88.850 90.830 ;
        RECT 91.105 90.740 92.235 90.830 ;
        RECT 106.480 90.915 110.565 91.615 ;
        RECT 106.480 89.770 107.180 90.915 ;
        RECT 109.435 90.740 110.565 90.915 ;
        RECT 87.890 88.580 89.020 89.750 ;
        RECT 106.220 88.600 107.350 89.770 ;
        RECT 88.165 86.995 88.865 88.580 ;
        RECT 90.425 86.995 91.555 87.370 ;
        RECT 88.165 86.295 91.555 86.995 ;
        RECT 106.495 87.135 107.195 88.600 ;
        RECT 108.755 87.135 109.885 87.370 ;
        RECT 106.495 86.435 109.885 87.135 ;
        RECT 90.425 86.200 91.555 86.295 ;
        RECT 108.755 86.200 109.885 86.435 ;
        RECT 90.780 85.220 91.480 86.200 ;
        RECT 92.500 85.220 93.630 85.945 ;
        RECT 90.780 84.775 93.630 85.220 ;
        RECT 109.110 85.360 109.810 86.200 ;
        RECT 110.830 85.360 111.960 85.945 ;
        RECT 109.110 84.775 111.960 85.360 ;
        RECT 90.780 84.520 93.415 84.775 ;
        RECT 109.110 84.660 111.745 84.775 ;
        RECT 92.715 84.000 93.415 84.520 ;
        RECT 111.045 84.000 111.745 84.660 ;
        RECT 65.200 83.175 66.330 83.630 ;
        RECT 74.245 83.380 75.375 83.780 ;
        RECT 63.820 82.875 66.330 83.175 ;
        RECT 52.275 76.635 53.755 76.935 ;
        RECT 52.275 76.400 53.005 76.635 ;
        RECT 45.720 73.900 46.850 74.335 ;
        RECT 53.455 74.200 53.755 76.635 ;
        RECT 54.705 74.210 55.835 74.310 ;
        RECT 63.820 74.210 64.120 82.875 ;
        RECT 65.200 82.460 66.330 82.875 ;
        RECT 72.695 83.080 75.375 83.380 ;
        RECT 65.200 74.210 66.330 74.455 ;
        RECT 54.705 74.200 66.330 74.210 ;
        RECT 53.455 73.910 66.330 74.200 ;
        RECT 53.455 73.900 55.835 73.910 ;
        RECT 45.720 73.780 53.755 73.900 ;
        RECT 44.755 73.600 53.755 73.780 ;
        RECT 44.755 73.480 46.850 73.600 ;
        RECT 45.720 73.165 46.850 73.480 ;
        RECT 54.705 73.140 55.835 73.900 ;
        RECT 65.200 73.285 66.330 73.910 ;
        RECT 72.695 73.690 72.995 83.080 ;
        RECT 74.245 82.610 75.375 83.080 ;
        RECT 92.500 82.830 93.630 84.000 ;
        RECT 110.830 82.830 111.960 84.000 ;
        RECT 92.580 82.085 93.280 82.830 ;
        RECT 94.770 82.085 95.900 82.460 ;
        RECT 92.580 81.385 95.900 82.085 ;
        RECT 94.770 81.290 95.900 81.385 ;
        RECT 97.925 82.105 99.055 82.460 ;
        RECT 110.910 82.105 111.610 82.830 ;
        RECT 113.100 82.105 114.230 82.460 ;
        RECT 97.925 81.405 114.230 82.105 ;
        RECT 97.925 81.290 99.055 81.405 ;
        RECT 94.985 80.965 95.685 81.290 ;
        RECT 98.150 80.965 98.850 81.290 ;
        RECT 94.985 80.265 98.850 80.965 ;
        RECT 96.150 78.220 97.280 78.415 ;
        RECT 94.410 77.520 97.280 78.220 ;
        RECT 94.410 76.690 95.110 77.520 ;
        RECT 96.150 77.245 97.280 77.520 ;
        RECT 94.195 76.465 95.325 76.690 ;
        RECT 93.180 75.765 95.325 76.465 ;
        RECT 93.180 75.255 93.880 75.765 ;
        RECT 94.195 75.520 95.325 75.765 ;
        RECT 90.835 75.125 93.885 75.255 ;
        RECT 90.835 74.555 94.295 75.125 ;
        RECT 73.840 73.690 74.970 74.155 ;
        RECT 72.695 73.390 74.970 73.690 ;
        RECT 90.835 73.620 91.535 74.555 ;
        RECT 93.165 73.955 94.295 74.555 ;
        RECT 72.695 72.840 72.995 73.390 ;
        RECT 73.840 72.985 74.970 73.390 ;
        RECT 90.815 73.385 91.945 73.620 ;
        RECT 50.425 72.540 72.995 72.840 ;
        RECT 87.665 72.685 91.945 73.385 ;
        RECT 50.425 66.700 50.725 72.540 ;
        RECT 58.380 70.275 58.680 72.540 ;
        RECT 87.665 71.480 88.365 72.685 ;
        RECT 90.815 72.450 91.945 72.685 ;
        RECT 87.600 70.310 88.730 71.480 ;
        RECT 58.195 69.505 58.925 70.275 ;
        RECT 87.665 68.615 88.365 70.310 ;
        RECT 90.135 68.615 91.265 69.080 ;
        RECT 87.665 67.915 91.265 68.615 ;
        RECT 90.135 67.910 91.265 67.915 ;
        RECT 51.315 66.700 52.445 67.135 ;
        RECT 50.425 66.400 52.445 66.700 ;
        RECT 47.755 59.960 48.485 60.240 ;
        RECT 50.425 59.960 50.725 66.400 ;
        RECT 51.315 65.965 52.445 66.400 ;
        RECT 90.490 66.840 91.190 67.910 ;
        RECT 92.210 66.840 93.340 67.655 ;
        RECT 90.490 66.485 93.340 66.840 ;
        RECT 90.490 66.140 93.125 66.485 ;
        RECT 92.425 65.710 93.125 66.140 ;
        RECT 92.210 64.540 93.340 65.710 ;
        RECT 92.290 63.705 92.990 64.540 ;
        RECT 94.480 63.705 95.610 64.170 ;
        RECT 92.290 63.005 95.610 63.705 ;
        RECT 94.480 63.000 95.610 63.005 ;
        RECT 97.635 63.470 98.765 64.170 ;
        RECT 103.255 63.470 103.955 81.405 ;
        RECT 113.100 81.290 114.230 81.405 ;
        RECT 116.255 81.290 117.385 82.460 ;
        RECT 113.445 80.985 114.145 81.290 ;
        RECT 116.470 80.985 117.170 81.290 ;
        RECT 113.445 80.285 117.170 80.985 ;
        RECT 114.750 77.975 115.880 78.170 ;
        RECT 113.060 77.275 115.880 77.975 ;
        RECT 113.060 76.445 113.760 77.275 ;
        RECT 114.750 77.000 115.880 77.275 ;
        RECT 112.845 76.220 113.975 76.445 ;
        RECT 111.805 75.520 113.975 76.220 ;
        RECT 111.805 75.010 112.505 75.520 ;
        RECT 112.845 75.275 113.975 75.520 ;
        RECT 109.465 74.880 112.515 75.010 ;
        RECT 109.465 74.310 112.945 74.880 ;
        RECT 109.465 73.375 110.165 74.310 ;
        RECT 111.805 74.295 112.945 74.310 ;
        RECT 111.815 73.710 112.945 74.295 ;
        RECT 109.465 73.140 110.595 73.375 ;
        RECT 106.295 72.440 110.595 73.140 ;
        RECT 106.295 71.250 106.995 72.440 ;
        RECT 109.465 72.205 110.595 72.440 ;
        RECT 106.250 70.080 107.380 71.250 ;
        RECT 106.295 68.600 106.995 70.080 ;
        RECT 108.785 68.600 109.915 68.835 ;
        RECT 106.295 67.900 109.915 68.600 ;
        RECT 108.785 67.665 109.915 67.900 ;
        RECT 109.140 66.825 109.840 67.665 ;
        RECT 110.860 66.825 111.990 67.410 ;
        RECT 109.140 66.240 111.990 66.825 ;
        RECT 109.140 66.125 111.775 66.240 ;
        RECT 111.075 65.465 111.775 66.125 ;
        RECT 110.860 64.295 111.990 65.465 ;
        RECT 110.940 63.470 111.640 64.295 ;
        RECT 113.130 63.470 114.260 63.925 ;
        RECT 97.635 63.000 114.260 63.470 ;
        RECT 94.695 62.585 95.395 63.000 ;
        RECT 97.850 62.770 114.260 63.000 ;
        RECT 97.850 62.585 98.560 62.770 ;
        RECT 94.695 61.885 98.560 62.585 ;
        RECT 102.365 62.105 103.065 62.770 ;
        RECT 113.130 62.755 114.260 62.770 ;
        RECT 116.285 62.755 117.415 63.925 ;
        RECT 113.345 62.350 114.045 62.755 ;
        RECT 116.510 62.350 117.210 62.755 ;
        RECT 102.365 61.365 103.140 62.105 ;
        RECT 113.345 61.650 117.210 62.350 ;
        RECT 102.420 61.325 103.140 61.365 ;
        RECT 51.315 59.960 52.445 60.445 ;
        RECT 47.755 59.660 52.445 59.960 ;
        RECT 47.755 59.470 48.485 59.660 ;
        RECT 51.315 59.275 52.445 59.660 ;
        RECT 105.130 60.075 109.800 60.105 ;
        RECT 105.130 59.405 112.400 60.075 ;
        RECT 105.130 56.660 105.830 59.405 ;
        RECT 108.720 59.375 112.400 59.405 ;
        RECT 108.720 58.290 109.420 59.375 ;
        RECT 111.700 58.290 112.400 59.375 ;
        RECT 108.485 57.120 109.615 58.290 ;
        RECT 111.485 57.120 112.615 58.290 ;
        RECT 106.235 56.660 107.365 56.880 ;
        RECT 72.770 55.315 73.890 56.495 ;
        RECT 103.935 55.960 107.365 56.660 ;
        RECT 103.935 54.770 104.635 55.960 ;
        RECT 106.235 55.710 107.365 55.960 ;
        RECT 105.900 54.770 107.030 55.205 ;
        RECT 103.935 54.470 107.030 54.770 ;
        RECT 51.315 53.345 52.445 53.780 ;
        RECT 50.415 53.045 52.445 53.345 ;
        RECT 50.415 46.865 50.715 53.045 ;
        RECT 51.315 52.610 52.445 53.045 ;
        RECT 61.330 50.720 62.460 51.890 ;
        RECT 72.770 51.565 73.890 52.745 ;
        RECT 103.935 51.730 104.635 54.470 ;
        RECT 105.900 54.035 107.030 54.470 ;
        RECT 103.935 51.150 104.700 51.730 ;
        RECT 105.900 51.150 107.030 51.585 ;
        RECT 103.935 51.030 107.030 51.150 ;
        RECT 59.815 49.395 60.945 50.565 ;
        RECT 61.745 50.005 62.045 50.720 ;
        RECT 60.355 47.850 60.655 49.395 ;
        RECT 61.330 48.835 62.460 50.005 ;
        RECT 72.865 49.835 73.995 51.005 ;
        RECT 103.995 50.850 107.030 51.030 ;
        RECT 61.745 48.180 62.045 48.835 ;
        RECT 73.330 48.435 73.630 49.835 ;
        RECT 61.330 47.850 62.460 48.180 ;
        RECT 60.355 47.550 62.460 47.850 ;
        RECT 51.315 46.955 52.445 47.155 ;
        RECT 60.355 46.955 60.655 47.550 ;
        RECT 61.330 47.010 62.460 47.550 ;
        RECT 72.805 47.265 73.935 48.435 ;
        RECT 51.315 46.865 60.655 46.955 ;
        RECT 50.415 46.655 60.655 46.865 ;
        RECT 50.415 46.565 52.445 46.655 ;
        RECT 51.315 45.985 52.445 46.565 ;
        RECT 61.745 46.305 62.045 47.010 ;
        RECT 61.330 45.135 62.460 46.305 ;
        RECT 73.330 45.930 73.630 47.265 ;
        RECT 103.995 45.995 104.695 50.850 ;
        RECT 105.900 50.415 107.030 50.850 ;
        RECT 105.900 47.600 107.030 47.835 ;
        RECT 105.555 46.665 107.030 47.600 ;
        RECT 105.555 45.995 106.255 46.665 ;
        RECT 106.575 45.995 107.705 46.230 ;
        RECT 61.745 44.485 62.045 45.135 ;
        RECT 72.915 44.760 74.045 45.930 ;
        RECT 103.995 45.295 107.705 45.995 ;
        RECT 61.330 43.315 62.460 44.485 ;
        RECT 73.330 43.320 73.630 44.760 ;
        RECT 61.745 42.745 62.045 43.315 ;
        RECT 61.330 41.575 62.460 42.745 ;
        RECT 72.915 42.150 74.045 43.320 ;
        RECT 36.850 40.490 38.490 40.520 ;
        RECT 39.240 40.490 40.370 40.925 ;
        RECT 48.050 40.500 49.180 40.935 ;
        RECT 61.745 40.910 62.045 41.575 ;
        RECT 36.850 40.190 40.370 40.490 ;
        RECT 36.850 34.020 37.150 40.190 ;
        RECT 39.240 39.755 40.370 40.190 ;
        RECT 45.875 40.200 49.180 40.500 ;
        RECT 38.890 34.020 40.020 34.220 ;
        RECT 36.850 33.720 40.020 34.020 ;
        RECT 36.850 27.800 37.150 33.720 ;
        RECT 38.890 33.050 40.020 33.720 ;
        RECT 45.875 33.805 46.175 40.200 ;
        RECT 48.050 39.765 49.180 40.200 ;
        RECT 61.330 39.740 62.460 40.910 ;
        RECT 73.330 40.835 73.630 42.150 ;
        RECT 97.110 41.730 98.240 42.220 ;
        RECT 105.555 41.730 106.255 45.295 ;
        RECT 106.575 45.060 107.705 45.295 ;
        RECT 108.985 43.570 110.115 44.740 ;
        RECT 111.715 43.610 112.845 44.780 ;
        RECT 109.230 41.730 109.930 43.570 ;
        RECT 111.930 41.730 112.630 43.610 ;
        RECT 97.110 41.050 112.630 41.730 ;
        RECT 97.325 41.030 112.630 41.050 ;
        RECT 72.915 39.665 74.045 40.835 ;
        RECT 73.330 38.950 73.630 39.665 ;
        RECT 73.000 38.180 73.730 38.950 ;
        RECT 58.890 36.265 60.020 36.700 ;
        RECT 72.730 36.265 73.860 37.060 ;
        RECT 56.075 35.965 73.860 36.265 ;
        RECT 48.035 33.860 49.165 34.230 ;
        RECT 56.075 33.860 56.375 35.965 ;
        RECT 58.890 35.530 60.020 35.965 ;
        RECT 72.730 35.890 73.860 35.965 ;
        RECT 45.875 33.795 47.060 33.805 ;
        RECT 48.035 33.795 56.375 33.860 ;
        RECT 45.875 33.560 56.375 33.795 ;
        RECT 45.875 33.495 49.165 33.560 ;
        RECT 38.890 27.800 40.020 28.105 ;
        RECT 36.850 27.500 40.020 27.800 ;
        RECT 36.850 21.275 37.150 27.500 ;
        RECT 38.890 26.935 40.020 27.500 ;
        RECT 45.875 27.770 46.175 33.495 ;
        RECT 48.035 33.060 49.165 33.495 ;
        RECT 57.705 33.220 58.425 33.345 ;
        RECT 58.890 33.220 60.020 33.655 ;
        RECT 57.705 32.920 60.020 33.220 ;
        RECT 57.705 32.565 58.425 32.920 ;
        RECT 58.890 32.485 60.020 32.920 ;
        RECT 48.070 27.770 49.200 28.135 ;
        RECT 45.875 27.470 49.200 27.770 ;
        RECT 37.900 21.275 39.030 21.710 ;
        RECT 36.850 21.190 39.030 21.275 ;
        RECT 45.875 21.190 46.175 27.470 ;
        RECT 46.805 27.450 47.105 27.470 ;
        RECT 48.070 26.965 49.200 27.470 ;
        RECT 48.025 21.190 49.155 21.730 ;
        RECT 36.850 20.975 49.155 21.190 ;
        RECT 37.900 20.890 49.155 20.975 ;
        RECT 37.900 20.540 39.030 20.890 ;
        RECT 48.025 20.560 49.155 20.890 ;
        RECT 97.110 19.425 98.240 19.860 ;
        RECT 102.040 19.425 124.495 35.925 ;
        RECT 97.110 19.125 124.495 19.425 ;
        RECT 97.110 18.690 98.240 19.125 ;
        RECT 102.040 13.475 124.495 19.125 ;
        RECT 134.190 4.545 135.360 4.550 ;
        RECT 154.745 4.545 155.915 4.550 ;
        RECT 112.215 4.205 113.385 4.210 ;
        RECT 112.210 3.085 113.390 4.205 ;
        RECT 134.185 3.425 135.365 4.545 ;
        RECT 154.740 3.425 155.920 4.545 ;
        RECT 134.190 3.420 135.360 3.425 ;
        RECT 154.745 3.420 155.915 3.425 ;
        RECT 112.215 3.080 113.385 3.085 ;
      LAYER via3 ;
        RECT 56.950 218.510 58.070 219.630 ;
        RECT 132.110 214.855 133.230 215.975 ;
        RECT 7.810 213.595 8.930 214.715 ;
        RECT 111.310 122.590 112.430 123.710 ;
        RECT 7.810 109.685 8.930 110.805 ;
        RECT 137.765 109.265 138.885 110.385 ;
        RECT 102.420 61.355 103.140 62.075 ;
        RECT 72.770 55.345 73.890 56.465 ;
        RECT 72.770 51.595 73.890 52.715 ;
        RECT 57.705 32.595 58.425 33.315 ;
        RECT 112.240 3.085 113.360 4.205 ;
        RECT 134.215 3.425 135.335 4.545 ;
        RECT 154.770 3.425 155.890 4.545 ;
      LAYER met4 ;
        RECT 3.980 225.045 3.990 225.750 ;
        RECT 7.660 225.045 7.670 225.750 ;
        RECT 11.340 225.045 11.350 225.750 ;
        RECT 15.020 225.045 15.030 225.750 ;
        RECT 18.700 225.045 18.710 225.750 ;
        RECT 22.380 225.045 22.390 225.750 ;
        RECT 26.060 225.045 26.070 225.750 ;
        RECT 29.740 225.045 29.750 225.750 ;
        RECT 33.420 225.045 33.430 225.750 ;
        RECT 37.100 225.045 37.110 225.750 ;
        RECT 40.780 225.045 40.790 225.750 ;
        RECT 44.460 225.045 44.470 225.750 ;
        RECT 48.140 225.045 48.150 225.750 ;
        RECT 51.820 225.045 51.830 225.750 ;
        RECT 55.500 225.045 55.510 225.750 ;
        RECT 59.180 225.045 59.190 225.750 ;
        RECT 62.860 225.045 62.870 225.750 ;
        RECT 66.540 225.045 66.550 225.750 ;
        RECT 70.220 225.045 70.230 225.750 ;
        RECT 73.900 225.045 73.910 225.750 ;
        RECT 77.580 225.045 77.590 225.750 ;
        RECT 81.260 225.045 81.270 225.750 ;
        RECT 84.940 225.045 84.950 225.750 ;
        RECT 88.620 225.045 88.630 225.750 ;
        RECT 3.480 224.760 3.990 225.045 ;
        RECT 4.290 224.760 7.670 225.045 ;
        RECT 7.970 224.760 11.350 225.045 ;
        RECT 11.650 224.760 15.030 225.045 ;
        RECT 15.330 224.760 18.710 225.045 ;
        RECT 19.010 224.760 22.390 225.045 ;
        RECT 22.690 224.760 26.070 225.045 ;
        RECT 26.370 224.760 29.750 225.045 ;
        RECT 30.050 224.760 33.430 225.045 ;
        RECT 33.730 224.760 37.110 225.045 ;
        RECT 37.410 224.760 40.790 225.045 ;
        RECT 41.090 224.760 44.470 225.045 ;
        RECT 44.770 224.760 48.150 225.045 ;
        RECT 48.450 224.760 51.830 225.045 ;
        RECT 52.130 224.760 55.510 225.045 ;
        RECT 55.810 224.760 59.190 225.045 ;
        RECT 59.490 224.760 62.870 225.045 ;
        RECT 63.170 224.760 66.550 225.045 ;
        RECT 66.850 224.760 70.230 225.045 ;
        RECT 70.530 224.760 73.910 225.045 ;
        RECT 74.210 224.760 77.590 225.045 ;
        RECT 77.890 224.760 81.270 225.045 ;
        RECT 81.570 224.760 84.950 225.045 ;
        RECT 85.250 224.760 88.630 225.045 ;
        RECT 92.300 224.760 92.310 225.750 ;
        RECT 95.980 224.760 95.990 225.750 ;
        RECT 99.660 224.760 99.670 225.750 ;
        RECT 103.340 224.760 103.350 225.750 ;
        RECT 107.020 224.760 107.030 225.750 ;
        RECT 110.700 224.760 110.710 225.750 ;
        RECT 114.380 224.760 114.390 225.750 ;
        RECT 118.060 224.760 118.070 225.750 ;
        RECT 121.740 224.760 121.750 225.750 ;
        RECT 125.420 224.760 125.430 225.750 ;
        RECT 129.100 224.760 129.110 225.750 ;
        RECT 132.780 224.760 132.790 225.750 ;
        RECT 136.460 224.760 136.470 225.750 ;
        RECT 140.140 224.760 140.150 225.750 ;
        RECT 143.820 224.760 143.830 225.750 ;
        RECT 147.500 224.760 147.510 225.750 ;
        RECT 151.180 224.760 151.190 225.750 ;
        RECT 154.860 224.760 154.870 225.750 ;
        RECT 158.540 224.760 158.550 225.750 ;
        RECT 3.480 224.750 88.920 224.760 ;
        RECT 92.300 224.750 92.600 224.760 ;
        RECT 95.980 224.750 96.280 224.760 ;
        RECT 99.660 224.750 99.960 224.760 ;
        RECT 103.340 224.750 103.640 224.760 ;
        RECT 107.020 224.750 107.320 224.760 ;
        RECT 110.700 224.750 111.000 224.760 ;
        RECT 114.380 224.750 114.680 224.760 ;
        RECT 118.060 224.750 118.360 224.760 ;
        RECT 121.740 224.750 122.040 224.760 ;
        RECT 125.420 224.750 125.720 224.760 ;
        RECT 129.100 224.750 129.400 224.760 ;
        RECT 132.780 224.750 133.080 224.760 ;
        RECT 136.460 224.750 136.760 224.760 ;
        RECT 140.140 224.750 140.440 224.760 ;
        RECT 143.820 224.750 144.120 224.760 ;
        RECT 147.500 224.750 147.800 224.760 ;
        RECT 151.180 224.750 151.480 224.760 ;
        RECT 154.860 224.750 155.160 224.760 ;
        RECT 158.540 224.750 158.840 224.760 ;
        RECT 3.480 224.745 88.760 224.750 ;
        RECT 3.480 214.655 5.480 224.745 ;
        RECT 56.945 219.570 58.075 219.635 ;
        RECT 15.015 218.570 58.075 219.570 ;
        RECT 7.805 214.655 8.935 214.720 ;
        RECT 3.480 213.655 8.935 214.655 ;
        RECT 3.480 110.745 5.480 213.655 ;
        RECT 7.805 213.590 8.935 213.655 ;
        RECT 7.805 110.745 8.935 110.810 ;
        RECT 3.480 109.745 8.935 110.745 ;
        RECT 1.990 0.000 2.000 0.990 ;
        RECT 3.480 0.205 5.480 109.745 ;
        RECT 7.805 109.680 8.935 109.745 ;
        RECT 15.015 2.665 16.015 218.570 ;
        RECT 56.945 218.505 58.075 218.570 ;
        RECT 132.105 215.915 133.235 215.980 ;
        RECT 158.345 215.915 160.345 224.140 ;
        RECT 132.105 214.915 160.345 215.915 ;
        RECT 132.105 214.850 133.235 214.915 ;
        RECT 111.305 123.650 112.435 123.715 ;
        RECT 20.490 122.650 112.435 123.650 ;
        RECT 20.490 4.560 21.490 122.650 ;
        RECT 111.305 122.585 112.435 122.650 ;
        RECT 137.760 110.325 138.890 110.390 ;
        RECT 158.345 110.325 160.345 214.915 ;
        RECT 137.760 109.325 160.345 110.325 ;
        RECT 137.760 109.260 138.890 109.325 ;
        RECT 102.415 61.350 103.145 62.080 ;
        RECT 72.765 55.340 73.895 56.470 ;
        RECT 73.180 53.435 73.480 55.340 ;
        RECT 59.380 53.135 73.480 53.435 ;
        RECT 59.380 44.910 59.680 53.135 ;
        RECT 73.180 52.720 73.480 53.135 ;
        RECT 72.765 51.590 73.895 52.720 ;
        RECT 57.760 44.890 59.680 44.910 ;
        RECT 56.745 44.610 59.680 44.890 ;
        RECT 56.745 44.590 58.060 44.610 ;
        RECT 56.745 33.105 57.045 44.590 ;
        RECT 102.430 35.785 103.130 61.350 ;
        RECT 57.700 33.105 58.430 33.320 ;
        RECT 56.745 32.805 58.430 33.105 ;
        RECT 57.700 32.590 58.430 32.805 ;
        RECT 102.180 13.615 124.355 35.785 ;
        RECT 20.490 3.560 91.090 4.560 ;
        RECT 15.015 1.665 69.035 2.665 ;
        RECT 68.035 1.000 69.035 1.665 ;
        RECT 24.070 0.000 24.080 0.990 ;
        RECT 46.150 0.000 46.160 0.990 ;
        RECT 68.035 0.485 68.240 1.000 ;
        RECT 68.840 0.485 69.035 1.000 ;
        RECT 90.090 1.000 91.090 3.560 ;
        RECT 112.235 3.080 113.365 4.210 ;
        RECT 134.210 3.420 135.340 4.550 ;
        RECT 154.765 4.485 155.895 4.550 ;
        RECT 154.765 3.485 157.395 4.485 ;
        RECT 154.765 3.420 155.895 3.485 ;
        RECT 90.090 0.550 90.320 1.000 ;
        RECT 90.920 0.550 91.090 1.000 ;
        RECT 112.300 1.000 113.300 3.080 ;
        RECT 112.300 0.755 112.400 1.000 ;
        RECT 113.000 0.755 113.300 1.000 ;
        RECT 134.275 1.000 135.275 3.420 ;
        RECT 68.230 0.000 68.240 0.485 ;
        RECT 90.310 0.000 90.320 0.550 ;
        RECT 112.390 0.000 112.400 0.755 ;
        RECT 134.275 0.450 134.480 1.000 ;
        RECT 135.080 0.450 135.275 1.000 ;
        RECT 156.395 1.000 157.395 3.485 ;
        RECT 156.395 0.460 156.560 1.000 ;
        RECT 157.160 0.460 157.395 1.000 ;
        RECT 134.470 0.000 134.480 0.450 ;
        RECT 156.550 0.000 156.560 0.460 ;
        RECT 158.345 0.255 160.345 109.325 ;
  END
END tt_um_Burrows_Katie
END LIBRARY

